//sin\cos�������ұ�
//�����ǽǶ�ֵ����2λ��1����0.25��
//���������ֵ����14λ
module lut_sin_cos(
    input             [10:0]       angle_div4,
    output reg signed [15:0]       sin_data,
    output reg signed [15:0]       cos_data
);

always@(angle_div4) begin
    case(angle_div4)
        11'd    0 , 11'd 720 : sin_data <= {16'd00000};
        11'd    1 , 11'd 719 : sin_data <= {16'd00071};
        11'd    2 , 11'd 718 : sin_data <= {16'd00143};
        11'd    3 , 11'd 717 : sin_data <= {16'd00214};
        11'd    4 , 11'd 716 : sin_data <= {16'd00286};
        11'd    5 , 11'd 715 : sin_data <= {16'd00357};
        11'd    6 , 11'd 714 : sin_data <= {16'd00429};
        11'd    7 , 11'd 713 : sin_data <= {16'd00500};
        11'd    8 , 11'd 712 : sin_data <= {16'd00572};
        11'd    9 , 11'd 711 : sin_data <= {16'd00643};
        11'd   10 , 11'd 710 : sin_data <= {16'd00715};
        11'd   11 , 11'd 709 : sin_data <= {16'd00786};
        11'd   12 , 11'd 708 : sin_data <= {16'd00857};
        11'd   13 , 11'd 707 : sin_data <= {16'd00929};
        11'd   14 , 11'd 706 : sin_data <= {16'd01000};
        11'd   15 , 11'd 705 : sin_data <= {16'd01072};
        11'd   16 , 11'd 704 : sin_data <= {16'd01143};
        11'd   17 , 11'd 703 : sin_data <= {16'd01214};
        11'd   18 , 11'd 702 : sin_data <= {16'd01285};
        11'd   19 , 11'd 701 : sin_data <= {16'd01357};
        11'd   20 , 11'd 700 : sin_data <= {16'd01428};
        11'd   21 , 11'd 699 : sin_data <= {16'd01499};
        11'd   22 , 11'd 698 : sin_data <= {16'd01570};
        11'd   23 , 11'd 697 : sin_data <= {16'd01641};
        11'd   24 , 11'd 696 : sin_data <= {16'd01713};
        11'd   25 , 11'd 695 : sin_data <= {16'd01784};
        11'd   26 , 11'd 694 : sin_data <= {16'd01855};
        11'd   27 , 11'd 693 : sin_data <= {16'd01926};
        11'd   28 , 11'd 692 : sin_data <= {16'd01997};
        11'd   29 , 11'd 691 : sin_data <= {16'd02068};
        11'd   30 , 11'd 690 : sin_data <= {16'd02139};
        11'd   31 , 11'd 689 : sin_data <= {16'd02209};
        11'd   32 , 11'd 688 : sin_data <= {16'd02280};
        11'd   33 , 11'd 687 : sin_data <= {16'd02351};
        11'd   34 , 11'd 686 : sin_data <= {16'd02422};
        11'd   35 , 11'd 685 : sin_data <= {16'd02492};
        11'd   36 , 11'd 684 : sin_data <= {16'd02563};
        11'd   37 , 11'd 683 : sin_data <= {16'd02634};
        11'd   38 , 11'd 682 : sin_data <= {16'd02704};
        11'd   39 , 11'd 681 : sin_data <= {16'd02775};
        11'd   40 , 11'd 680 : sin_data <= {16'd02845};
        11'd   41 , 11'd 679 : sin_data <= {16'd02915};
        11'd   42 , 11'd 678 : sin_data <= {16'd02986};
        11'd   43 , 11'd 677 : sin_data <= {16'd03056};
        11'd   44 , 11'd 676 : sin_data <= {16'd03126};
        11'd   45 , 11'd 675 : sin_data <= {16'd03196};
        11'd   46 , 11'd 674 : sin_data <= {16'd03266};
        11'd   47 , 11'd 673 : sin_data <= {16'd03336};
        11'd   48 , 11'd 672 : sin_data <= {16'd03406};
        11'd   49 , 11'd 671 : sin_data <= {16'd03476};
        11'd   50 , 11'd 670 : sin_data <= {16'd03546};
        11'd   51 , 11'd 669 : sin_data <= {16'd03616};
        11'd   52 , 11'd 668 : sin_data <= {16'd03686};
        11'd   53 , 11'd 667 : sin_data <= {16'd03755};
        11'd   54 , 11'd 666 : sin_data <= {16'd03825};
        11'd   55 , 11'd 665 : sin_data <= {16'd03894};
        11'd   56 , 11'd 664 : sin_data <= {16'd03964};
        11'd   57 , 11'd 663 : sin_data <= {16'd04033};
        11'd   58 , 11'd 662 : sin_data <= {16'd04102};
        11'd   59 , 11'd 661 : sin_data <= {16'd04171};
        11'd   60 , 11'd 660 : sin_data <= {16'd04240};
        11'd   61 , 11'd 659 : sin_data <= {16'd04310};
        11'd   62 , 11'd 658 : sin_data <= {16'd04378};
        11'd   63 , 11'd 657 : sin_data <= {16'd04447};
        11'd   64 , 11'd 656 : sin_data <= {16'd04516};
        11'd   65 , 11'd 655 : sin_data <= {16'd04585};
        11'd   66 , 11'd 654 : sin_data <= {16'd04653};
        11'd   67 , 11'd 653 : sin_data <= {16'd04722};
        11'd   68 , 11'd 652 : sin_data <= {16'd04790};
        11'd   69 , 11'd 651 : sin_data <= {16'd04859};
        11'd   70 , 11'd 650 : sin_data <= {16'd04927};
        11'd   71 , 11'd 649 : sin_data <= {16'd04995};
        11'd   72 , 11'd 648 : sin_data <= {16'd05063};
        11'd   73 , 11'd 647 : sin_data <= {16'd05131};
        11'd   74 , 11'd 646 : sin_data <= {16'd05199};
        11'd   75 , 11'd 645 : sin_data <= {16'd05266};
        11'd   76 , 11'd 644 : sin_data <= {16'd05334};
        11'd   77 , 11'd 643 : sin_data <= {16'd05402};
        11'd   78 , 11'd 642 : sin_data <= {16'd05469};
        11'd   79 , 11'd 641 : sin_data <= {16'd05536};
        11'd   80 , 11'd 640 : sin_data <= {16'd05604};
        11'd   81 , 11'd 639 : sin_data <= {16'd05671};
        11'd   82 , 11'd 638 : sin_data <= {16'd05738};
        11'd   83 , 11'd 637 : sin_data <= {16'd05805};
        11'd   84 , 11'd 636 : sin_data <= {16'd05872};
        11'd   85 , 11'd 635 : sin_data <= {16'd05938};
        11'd   86 , 11'd 634 : sin_data <= {16'd06005};
        11'd   87 , 11'd 633 : sin_data <= {16'd06071};
        11'd   88 , 11'd 632 : sin_data <= {16'd06138};
        11'd   89 , 11'd 631 : sin_data <= {16'd06204};
        11'd   90 , 11'd 630 : sin_data <= {16'd06270};
        11'd   91 , 11'd 629 : sin_data <= {16'd06336};
        11'd   92 , 11'd 628 : sin_data <= {16'd06402};
        11'd   93 , 11'd 627 : sin_data <= {16'd06467};
        11'd   94 , 11'd 626 : sin_data <= {16'd06533};
        11'd   95 , 11'd 625 : sin_data <= {16'd06599};
        11'd   96 , 11'd 624 : sin_data <= {16'd06664};
        11'd   97 , 11'd 623 : sin_data <= {16'd06729};
        11'd   98 , 11'd 622 : sin_data <= {16'd06794};
        11'd   99 , 11'd 621 : sin_data <= {16'd06859};
        11'd  100 , 11'd 620 : sin_data <= {16'd06924};
        11'd  101 , 11'd 619 : sin_data <= {16'd06989};
        11'd  102 , 11'd 618 : sin_data <= {16'd07053};
        11'd  103 , 11'd 617 : sin_data <= {16'd07118};
        11'd  104 , 11'd 616 : sin_data <= {16'd07182};
        11'd  105 , 11'd 615 : sin_data <= {16'd07246};
        11'd  106 , 11'd 614 : sin_data <= {16'd07311};
        11'd  107 , 11'd 613 : sin_data <= {16'd07374};
        11'd  108 , 11'd 612 : sin_data <= {16'd07438};
        11'd  109 , 11'd 611 : sin_data <= {16'd07502};
        11'd  110 , 11'd 610 : sin_data <= {16'd07565};
        11'd  111 , 11'd 609 : sin_data <= {16'd07629};
        11'd  112 , 11'd 608 : sin_data <= {16'd07692};
        11'd  113 , 11'd 607 : sin_data <= {16'd07755};
        11'd  114 , 11'd 606 : sin_data <= {16'd07818};
        11'd  115 , 11'd 605 : sin_data <= {16'd07881};
        11'd  116 , 11'd 604 : sin_data <= {16'd07943};
        11'd  117 , 11'd 603 : sin_data <= {16'd08006};
        11'd  118 , 11'd 602 : sin_data <= {16'd08068};
        11'd  119 , 11'd 601 : sin_data <= {16'd08130};
        11'd  120 , 11'd 600 : sin_data <= {16'd08192};
        11'd  121 , 11'd 599 : sin_data <= {16'd08254};
        11'd  122 , 11'd 598 : sin_data <= {16'd08316};
        11'd  123 , 11'd 597 : sin_data <= {16'd08377};
        11'd  124 , 11'd 596 : sin_data <= {16'd08438};
        11'd  125 , 11'd 595 : sin_data <= {16'd08500};
        11'd  126 , 11'd 594 : sin_data <= {16'd08561};
        11'd  127 , 11'd 593 : sin_data <= {16'd08621};
        11'd  128 , 11'd 592 : sin_data <= {16'd08682};
        11'd  129 , 11'd 591 : sin_data <= {16'd08743};
        11'd  130 , 11'd 590 : sin_data <= {16'd08803};
        11'd  131 , 11'd 589 : sin_data <= {16'd08863};
        11'd  132 , 11'd 588 : sin_data <= {16'd08923};
        11'd  133 , 11'd 587 : sin_data <= {16'd08983};
        11'd  134 , 11'd 586 : sin_data <= {16'd09043};
        11'd  135 , 11'd 585 : sin_data <= {16'd09102};
        11'd  136 , 11'd 584 : sin_data <= {16'd09162};
        11'd  137 , 11'd 583 : sin_data <= {16'd09221};
        11'd  138 , 11'd 582 : sin_data <= {16'd09280};
        11'd  139 , 11'd 581 : sin_data <= {16'd09339};
        11'd  140 , 11'd 580 : sin_data <= {16'd09397};
        11'd  141 , 11'd 579 : sin_data <= {16'd09456};
        11'd  142 , 11'd 578 : sin_data <= {16'd09514};
        11'd  143 , 11'd 577 : sin_data <= {16'd09572};
        11'd  144 , 11'd 576 : sin_data <= {16'd09630};
        11'd  145 , 11'd 575 : sin_data <= {16'd09688};
        11'd  146 , 11'd 574 : sin_data <= {16'd09746};
        11'd  147 , 11'd 573 : sin_data <= {16'd09803};
        11'd  148 , 11'd 572 : sin_data <= {16'd09860};
        11'd  149 , 11'd 571 : sin_data <= {16'd09917};
        11'd  150 , 11'd 570 : sin_data <= {16'd09974};
        11'd  151 , 11'd 569 : sin_data <= {16'd10031};
        11'd  152 , 11'd 568 : sin_data <= {16'd10087};
        11'd  153 , 11'd 567 : sin_data <= {16'd10143};
        11'd  154 , 11'd 566 : sin_data <= {16'd10199};
        11'd  155 , 11'd 565 : sin_data <= {16'd10255};
        11'd  156 , 11'd 564 : sin_data <= {16'd10311};
        11'd  157 , 11'd 563 : sin_data <= {16'd10366};
        11'd  158 , 11'd 562 : sin_data <= {16'd10422};
        11'd  159 , 11'd 561 : sin_data <= {16'd10477};
        11'd  160 , 11'd 560 : sin_data <= {16'd10531};
        11'd  161 , 11'd 559 : sin_data <= {16'd10586};
        11'd  162 , 11'd 558 : sin_data <= {16'd10641};
        11'd  163 , 11'd 557 : sin_data <= {16'd10695};
        11'd  164 , 11'd 556 : sin_data <= {16'd10749};
        11'd  165 , 11'd 555 : sin_data <= {16'd10803};
        11'd  166 , 11'd 554 : sin_data <= {16'd10856};
        11'd  167 , 11'd 553 : sin_data <= {16'd10910};
        11'd  168 , 11'd 552 : sin_data <= {16'd10963};
        11'd  169 , 11'd 551 : sin_data <= {16'd11016};
        11'd  170 , 11'd 550 : sin_data <= {16'd11069};
        11'd  171 , 11'd 549 : sin_data <= {16'd11121};
        11'd  172 , 11'd 548 : sin_data <= {16'd11174};
        11'd  173 , 11'd 547 : sin_data <= {16'd11226};
        11'd  174 , 11'd 546 : sin_data <= {16'd11278};
        11'd  175 , 11'd 545 : sin_data <= {16'd11330};
        11'd  176 , 11'd 544 : sin_data <= {16'd11381};
        11'd  177 , 11'd 543 : sin_data <= {16'd11433};
        11'd  178 , 11'd 542 : sin_data <= {16'd11484};
        11'd  179 , 11'd 541 : sin_data <= {16'd11535};
        11'd  180 , 11'd 540 : sin_data <= {16'd11585};
        11'd  181 , 11'd 539 : sin_data <= {16'd11636};
        11'd  182 , 11'd 538 : sin_data <= {16'd11686};
        11'd  183 , 11'd 537 : sin_data <= {16'd11736};
        11'd  184 , 11'd 536 : sin_data <= {16'd11786};
        11'd  185 , 11'd 535 : sin_data <= {16'd11835};
        11'd  186 , 11'd 534 : sin_data <= {16'd11885};
        11'd  187 , 11'd 533 : sin_data <= {16'd11934};
        11'd  188 , 11'd 532 : sin_data <= {16'd11982};
        11'd  189 , 11'd 531 : sin_data <= {16'd12031};
        11'd  190 , 11'd 530 : sin_data <= {16'd12080};
        11'd  191 , 11'd 529 : sin_data <= {16'd12128};
        11'd  192 , 11'd 528 : sin_data <= {16'd12176};
        11'd  193 , 11'd 527 : sin_data <= {16'd12223};
        11'd  194 , 11'd 526 : sin_data <= {16'd12271};
        11'd  195 , 11'd 525 : sin_data <= {16'd12318};
        11'd  196 , 11'd 524 : sin_data <= {16'd12365};
        11'd  197 , 11'd 523 : sin_data <= {16'd12412};
        11'd  198 , 11'd 522 : sin_data <= {16'd12458};
        11'd  199 , 11'd 521 : sin_data <= {16'd12505};
        11'd  200 , 11'd 520 : sin_data <= {16'd12551};
        11'd  201 , 11'd 519 : sin_data <= {16'd12597};
        11'd  202 , 11'd 518 : sin_data <= {16'd12642};
        11'd  203 , 11'd 517 : sin_data <= {16'd12688};
        11'd  204 , 11'd 516 : sin_data <= {16'd12733};
        11'd  205 , 11'd 515 : sin_data <= {16'd12778};
        11'd  206 , 11'd 514 : sin_data <= {16'd12822};
        11'd  207 , 11'd 513 : sin_data <= {16'd12867};
        11'd  208 , 11'd 512 : sin_data <= {16'd12911};
        11'd  209 , 11'd 511 : sin_data <= {16'd12955};
        11'd  210 , 11'd 510 : sin_data <= {16'd12998};
        11'd  211 , 11'd 509 : sin_data <= {16'd13042};
        11'd  212 , 11'd 508 : sin_data <= {16'd13085};
        11'd  213 , 11'd 507 : sin_data <= {16'd13128};
        11'd  214 , 11'd 506 : sin_data <= {16'd13170};
        11'd  215 , 11'd 505 : sin_data <= {16'd13213};
        11'd  216 , 11'd 504 : sin_data <= {16'd13255};
        11'd  217 , 11'd 503 : sin_data <= {16'd13297};
        11'd  218 , 11'd 502 : sin_data <= {16'd13338};
        11'd  219 , 11'd 501 : sin_data <= {16'd13380};
        11'd  220 , 11'd 500 : sin_data <= {16'd13421};
        11'd  221 , 11'd 499 : sin_data <= {16'd13462};
        11'd  222 , 11'd 498 : sin_data <= {16'd13502};
        11'd  223 , 11'd 497 : sin_data <= {16'd13543};
        11'd  224 , 11'd 496 : sin_data <= {16'd13583};
        11'd  225 , 11'd 495 : sin_data <= {16'd13623};
        11'd  226 , 11'd 494 : sin_data <= {16'd13662};
        11'd  227 , 11'd 493 : sin_data <= {16'd13702};
        11'd  228 , 11'd 492 : sin_data <= {16'd13741};
        11'd  229 , 11'd 491 : sin_data <= {16'd13780};
        11'd  230 , 11'd 490 : sin_data <= {16'd13818};
        11'd  231 , 11'd 489 : sin_data <= {16'd13856};
        11'd  232 , 11'd 488 : sin_data <= {16'd13894};
        11'd  233 , 11'd 487 : sin_data <= {16'd13932};
        11'd  234 , 11'd 486 : sin_data <= {16'd13970};
        11'd  235 , 11'd 485 : sin_data <= {16'd14007};
        11'd  236 , 11'd 484 : sin_data <= {16'd14044};
        11'd  237 , 11'd 483 : sin_data <= {16'd14081};
        11'd  238 , 11'd 482 : sin_data <= {16'd14117};
        11'd  239 , 11'd 481 : sin_data <= {16'd14153};
        11'd  240 , 11'd 480 : sin_data <= {16'd14189};
        11'd  241 , 11'd 479 : sin_data <= {16'd14225};
        11'd  242 , 11'd 478 : sin_data <= {16'd14260};
        11'd  243 , 11'd 477 : sin_data <= {16'd14295};
        11'd  244 , 11'd 476 : sin_data <= {16'd14330};
        11'd  245 , 11'd 475 : sin_data <= {16'd14364};
        11'd  246 , 11'd 474 : sin_data <= {16'd14399};
        11'd  247 , 11'd 473 : sin_data <= {16'd14433};
        11'd  248 , 11'd 472 : sin_data <= {16'd14466};
        11'd  249 , 11'd 471 : sin_data <= {16'd14500};
        11'd  250 , 11'd 470 : sin_data <= {16'd14533};
        11'd  251 , 11'd 469 : sin_data <= {16'd14566};
        11'd  252 , 11'd 468 : sin_data <= {16'd14598};
        11'd  253 , 11'd 467 : sin_data <= {16'd14631};
        11'd  254 , 11'd 466 : sin_data <= {16'd14663};
        11'd  255 , 11'd 465 : sin_data <= {16'd14694};
        11'd  256 , 11'd 464 : sin_data <= {16'd14726};
        11'd  257 , 11'd 463 : sin_data <= {16'd14757};
        11'd  258 , 11'd 462 : sin_data <= {16'd14788};
        11'd  259 , 11'd 461 : sin_data <= {16'd14819};
        11'd  260 , 11'd 460 : sin_data <= {16'd14849};
        11'd  261 , 11'd 459 : sin_data <= {16'd14879};
        11'd  262 , 11'd 458 : sin_data <= {16'd14909};
        11'd  263 , 11'd 457 : sin_data <= {16'd14938};
        11'd  264 , 11'd 456 : sin_data <= {16'd14968};
        11'd  265 , 11'd 455 : sin_data <= {16'd14996};
        11'd  266 , 11'd 454 : sin_data <= {16'd15025};
        11'd  267 , 11'd 453 : sin_data <= {16'd15053};
        11'd  268 , 11'd 452 : sin_data <= {16'd15082};
        11'd  269 , 11'd 451 : sin_data <= {16'd15109};
        11'd  270 , 11'd 450 : sin_data <= {16'd15137};
        11'd  271 , 11'd 449 : sin_data <= {16'd15164};
        11'd  272 , 11'd 448 : sin_data <= {16'd15191};
        11'd  273 , 11'd 447 : sin_data <= {16'd15218};
        11'd  274 , 11'd 446 : sin_data <= {16'd15244};
        11'd  275 , 11'd 445 : sin_data <= {16'd15270};
        11'd  276 , 11'd 444 : sin_data <= {16'd15296};
        11'd  277 , 11'd 443 : sin_data <= {16'd15321};
        11'd  278 , 11'd 442 : sin_data <= {16'd15346};
        11'd  279 , 11'd 441 : sin_data <= {16'd15371};
        11'd  280 , 11'd 440 : sin_data <= {16'd15396};
        11'd  281 , 11'd 439 : sin_data <= {16'd15420};
        11'd  282 , 11'd 438 : sin_data <= {16'd15444};
        11'd  283 , 11'd 437 : sin_data <= {16'd15468};
        11'd  284 , 11'd 436 : sin_data <= {16'd15491};
        11'd  285 , 11'd 435 : sin_data <= {16'd15515};
        11'd  286 , 11'd 434 : sin_data <= {16'd15537};
        11'd  287 , 11'd 433 : sin_data <= {16'd15560};
        11'd  288 , 11'd 432 : sin_data <= {16'd15582};
        11'd  289 , 11'd 431 : sin_data <= {16'd15604};
        11'd  290 , 11'd 430 : sin_data <= {16'd15626};
        11'd  291 , 11'd 429 : sin_data <= {16'd15647};
        11'd  292 , 11'd 428 : sin_data <= {16'd15668};
        11'd  293 , 11'd 427 : sin_data <= {16'd15689};
        11'd  294 , 11'd 426 : sin_data <= {16'd15709};
        11'd  295 , 11'd 425 : sin_data <= {16'd15729};
        11'd  296 , 11'd 424 : sin_data <= {16'd15749};
        11'd  297 , 11'd 423 : sin_data <= {16'd15769};
        11'd  298 , 11'd 422 : sin_data <= {16'd15788};
        11'd  299 , 11'd 421 : sin_data <= {16'd15807};
        11'd  300 , 11'd 420 : sin_data <= {16'd15826};
        11'd  301 , 11'd 419 : sin_data <= {16'd15844};
        11'd  302 , 11'd 418 : sin_data <= {16'd15862};
        11'd  303 , 11'd 417 : sin_data <= {16'd15880};
        11'd  304 , 11'd 416 : sin_data <= {16'd15897};
        11'd  305 , 11'd 415 : sin_data <= {16'd15914};
        11'd  306 , 11'd 414 : sin_data <= {16'd15931};
        11'd  307 , 11'd 413 : sin_data <= {16'd15948};
        11'd  308 , 11'd 412 : sin_data <= {16'd15964};
        11'd  309 , 11'd 411 : sin_data <= {16'd15980};
        11'd  310 , 11'd 410 : sin_data <= {16'd15996};
        11'd  311 , 11'd 409 : sin_data <= {16'd16011};
        11'd  312 , 11'd 408 : sin_data <= {16'd16026};
        11'd  313 , 11'd 407 : sin_data <= {16'd16041};
        11'd  314 , 11'd 406 : sin_data <= {16'd16055};
        11'd  315 , 11'd 405 : sin_data <= {16'd16069};
        11'd  316 , 11'd 404 : sin_data <= {16'd16083};
        11'd  317 , 11'd 403 : sin_data <= {16'd16096};
        11'd  318 , 11'd 402 : sin_data <= {16'd16110};
        11'd  319 , 11'd 401 : sin_data <= {16'd16123};
        11'd  320 , 11'd 400 : sin_data <= {16'd16135};
        11'd  321 , 11'd 399 : sin_data <= {16'd16147};
        11'd  322 , 11'd 398 : sin_data <= {16'd16159};
        11'd  323 , 11'd 397 : sin_data <= {16'd16171};
        11'd  324 , 11'd 396 : sin_data <= {16'd16182};
        11'd  325 , 11'd 395 : sin_data <= {16'd16193};
        11'd  326 , 11'd 394 : sin_data <= {16'd16204};
        11'd  327 , 11'd 393 : sin_data <= {16'd16214};
        11'd  328 , 11'd 392 : sin_data <= {16'd16225};
        11'd  329 , 11'd 391 : sin_data <= {16'd16234};
        11'd  330 , 11'd 390 : sin_data <= {16'd16244};
        11'd  331 , 11'd 389 : sin_data <= {16'd16253};
        11'd  332 , 11'd 388 : sin_data <= {16'd16262};
        11'd  333 , 11'd 387 : sin_data <= {16'd16270};
        11'd  334 , 11'd 386 : sin_data <= {16'd16279};
        11'd  335 , 11'd 385 : sin_data <= {16'd16287};
        11'd  336 , 11'd 384 : sin_data <= {16'd16294};
        11'd  337 , 11'd 383 : sin_data <= {16'd16302};
        11'd  338 , 11'd 382 : sin_data <= {16'd16309};
        11'd  339 , 11'd 381 : sin_data <= {16'd16315};
        11'd  340 , 11'd 380 : sin_data <= {16'd16322};
        11'd  341 , 11'd 379 : sin_data <= {16'd16328};
        11'd  342 , 11'd 378 : sin_data <= {16'd16333};
        11'd  343 , 11'd 377 : sin_data <= {16'd16339};
        11'd  344 , 11'd 376 : sin_data <= {16'd16344};
        11'd  345 , 11'd 375 : sin_data <= {16'd16349};
        11'd  346 , 11'd 374 : sin_data <= {16'd16353};
        11'd  347 , 11'd 373 : sin_data <= {16'd16358};
        11'd  348 , 11'd 372 : sin_data <= {16'd16362};
        11'd  349 , 11'd 371 : sin_data <= {16'd16365};
        11'd  350 , 11'd 370 : sin_data <= {16'd16368};
        11'd  351 , 11'd 369 : sin_data <= {16'd16371};
        11'd  352 , 11'd 368 : sin_data <= {16'd16374};
        11'd  353 , 11'd 367 : sin_data <= {16'd16376};
        11'd  354 , 11'd 366 : sin_data <= {16'd16378};
        11'd  355 , 11'd 365 : sin_data <= {16'd16380};
        11'd  356 , 11'd 364 : sin_data <= {16'd16382};
        11'd  357 , 11'd 363 : sin_data <= {16'd16383};
        11'd  358 , 11'd 362 : sin_data <= {16'd16383};
        11'd  359 , 11'd 361 : sin_data <= {16'd16384};
        11'd  360            : sin_data <= {16'd16384};
        



                    11'd 1440 : sin_data <= {-16'd00000};    
        11'd  721 , 11'd 1439 : sin_data <= {-16'd00071};
        11'd  722 , 11'd 1438 : sin_data <= {-16'd00143};
        11'd  723 , 11'd 1437 : sin_data <= {-16'd00214};
        11'd  724 , 11'd 1436 : sin_data <= {-16'd00286};
        11'd  725 , 11'd 1435 : sin_data <= {-16'd00357};
        11'd  726 , 11'd 1434 : sin_data <= {-16'd00429};
        11'd  727 , 11'd 1433 : sin_data <= {-16'd00500};
        11'd  728 , 11'd 1432 : sin_data <= {-16'd00572};
        11'd  729 , 11'd 1431 : sin_data <= {-16'd00643};
        11'd  730 , 11'd 1430 : sin_data <= {-16'd00715};
        11'd  731 , 11'd 1429 : sin_data <= {-16'd00786};
        11'd  732 , 11'd 1428 : sin_data <= {-16'd00857};
        11'd  733 , 11'd 1427 : sin_data <= {-16'd00929};
        11'd  734 , 11'd 1426 : sin_data <= {-16'd01000};
        11'd  735 , 11'd 1425 : sin_data <= {-16'd01072};
        11'd  736 , 11'd 1424 : sin_data <= {-16'd01143};
        11'd  737 , 11'd 1423 : sin_data <= {-16'd01214};
        11'd  738 , 11'd 1422 : sin_data <= {-16'd01285};
        11'd  739 , 11'd 1421 : sin_data <= {-16'd01357};
        11'd  740 , 11'd 1420 : sin_data <= {-16'd01428};
        11'd  741 , 11'd 1419 : sin_data <= {-16'd01499};
        11'd  742 , 11'd 1418 : sin_data <= {-16'd01570};
        11'd  743 , 11'd 1417 : sin_data <= {-16'd01641};
        11'd  744 , 11'd 1416 : sin_data <= {-16'd01713};
        11'd  745 , 11'd 1415 : sin_data <= {-16'd01784};
        11'd  746 , 11'd 1414 : sin_data <= {-16'd01855};
        11'd  747 , 11'd 1413 : sin_data <= {-16'd01926};
        11'd  748 , 11'd 1412 : sin_data <= {-16'd01997};
        11'd  749 , 11'd 1411 : sin_data <= {-16'd02068};
        11'd  750 , 11'd 1410 : sin_data <= {-16'd02139};
        11'd  751 , 11'd 1409 : sin_data <= {-16'd02209};
        11'd  752 , 11'd 1408 : sin_data <= {-16'd02280};
        11'd  753 , 11'd 1407 : sin_data <= {-16'd02351};
        11'd  754 , 11'd 1406 : sin_data <= {-16'd02422};
        11'd  755 , 11'd 1405 : sin_data <= {-16'd02492};
        11'd  756 , 11'd 1404 : sin_data <= {-16'd02563};
        11'd  757 , 11'd 1403 : sin_data <= {-16'd02634};
        11'd  758 , 11'd 1402 : sin_data <= {-16'd02704};
        11'd  759 , 11'd 1401 : sin_data <= {-16'd02775};
        11'd  760 , 11'd 1400 : sin_data <= {-16'd02845};
        11'd  761 , 11'd 1399 : sin_data <= {-16'd02915};
        11'd  762 , 11'd 1398 : sin_data <= {-16'd02986};
        11'd  763 , 11'd 1397 : sin_data <= {-16'd03056};
        11'd  764 , 11'd 1396 : sin_data <= {-16'd03126};
        11'd  765 , 11'd 1395 : sin_data <= {-16'd03196};
        11'd  766 , 11'd 1394 : sin_data <= {-16'd03266};
        11'd  767 , 11'd 1393 : sin_data <= {-16'd03336};
        11'd  768 , 11'd 1392 : sin_data <= {-16'd03406};
        11'd  769 , 11'd 1391 : sin_data <= {-16'd03476};
        11'd  770 , 11'd 1390 : sin_data <= {-16'd03546};
        11'd  771 , 11'd 1389 : sin_data <= {-16'd03616};
        11'd  772 , 11'd 1388 : sin_data <= {-16'd03686};
        11'd  773 , 11'd 1387 : sin_data <= {-16'd03755};
        11'd  774 , 11'd 1386 : sin_data <= {-16'd03825};
        11'd  775 , 11'd 1385 : sin_data <= {-16'd03894};
        11'd  776 , 11'd 1384 : sin_data <= {-16'd03964};
        11'd  777 , 11'd 1383 : sin_data <= {-16'd04033};
        11'd  778 , 11'd 1382 : sin_data <= {-16'd04102};
        11'd  779 , 11'd 1381 : sin_data <= {-16'd04171};
        11'd  780 , 11'd 1380 : sin_data <= {-16'd04240};
        11'd  781 , 11'd 1379 : sin_data <= {-16'd04310};
        11'd  782 , 11'd 1378 : sin_data <= {-16'd04378};
        11'd  783 , 11'd 1377 : sin_data <= {-16'd04447};
        11'd  784 , 11'd 1376 : sin_data <= {-16'd04516};
        11'd  785 , 11'd 1375 : sin_data <= {-16'd04585};
        11'd  786 , 11'd 1374 : sin_data <= {-16'd04653};
        11'd  787 , 11'd 1373 : sin_data <= {-16'd04722};
        11'd  788 , 11'd 1372 : sin_data <= {-16'd04790};
        11'd  789 , 11'd 1371 : sin_data <= {-16'd04859};
        11'd  790 , 11'd 1370 : sin_data <= {-16'd04927};
        11'd  791 , 11'd 1369 : sin_data <= {-16'd04995};
        11'd  792 , 11'd 1368 : sin_data <= {-16'd05063};
        11'd  793 , 11'd 1367 : sin_data <= {-16'd05131};
        11'd  794 , 11'd 1366 : sin_data <= {-16'd05199};
        11'd  795 , 11'd 1365 : sin_data <= {-16'd05266};
        11'd  796 , 11'd 1364 : sin_data <= {-16'd05334};
        11'd  797 , 11'd 1363 : sin_data <= {-16'd05402};
        11'd  798 , 11'd 1362 : sin_data <= {-16'd05469};
        11'd  799 , 11'd 1361 : sin_data <= {-16'd05536};
        11'd  800 , 11'd 1360 : sin_data <= {-16'd05604};
        11'd  801 , 11'd 1359 : sin_data <= {-16'd05671};
        11'd  802 , 11'd 1358 : sin_data <= {-16'd05738};
        11'd  803 , 11'd 1357 : sin_data <= {-16'd05805};
        11'd  804 , 11'd 1356 : sin_data <= {-16'd05872};
        11'd  805 , 11'd 1355 : sin_data <= {-16'd05938};
        11'd  806 , 11'd 1354 : sin_data <= {-16'd06005};
        11'd  807 , 11'd 1353 : sin_data <= {-16'd06071};
        11'd  808 , 11'd 1352 : sin_data <= {-16'd06138};
        11'd  809 , 11'd 1351 : sin_data <= {-16'd06204};
        11'd  810 , 11'd 1350 : sin_data <= {-16'd06270};
        11'd  811 , 11'd 1349 : sin_data <= {-16'd06336};
        11'd  812 , 11'd 1348 : sin_data <= {-16'd06402};
        11'd  813 , 11'd 1347 : sin_data <= {-16'd06467};
        11'd  814 , 11'd 1346 : sin_data <= {-16'd06533};
        11'd  815 , 11'd 1345 : sin_data <= {-16'd06599};
        11'd  816 , 11'd 1344 : sin_data <= {-16'd06664};
        11'd  817 , 11'd 1343 : sin_data <= {-16'd06729};
        11'd  818 , 11'd 1342 : sin_data <= {-16'd06794};
        11'd  819 , 11'd 1341 : sin_data <= {-16'd06859};
        11'd  820 , 11'd 1340 : sin_data <= {-16'd06924};
        11'd  821 , 11'd 1339 : sin_data <= {-16'd06989};
        11'd  822 , 11'd 1338 : sin_data <= {-16'd07053};
        11'd  823 , 11'd 1337 : sin_data <= {-16'd07118};
        11'd  824 , 11'd 1336 : sin_data <= {-16'd07182};
        11'd  825 , 11'd 1335 : sin_data <= {-16'd07246};
        11'd  826 , 11'd 1334 : sin_data <= {-16'd07311};
        11'd  827 , 11'd 1333 : sin_data <= {-16'd07374};
        11'd  828 , 11'd 1332 : sin_data <= {-16'd07438};
        11'd  829 , 11'd 1331 : sin_data <= {-16'd07502};
        11'd  830 , 11'd 1330 : sin_data <= {-16'd07565};
        11'd  831 , 11'd 1329 : sin_data <= {-16'd07629};
        11'd  832 , 11'd 1328 : sin_data <= {-16'd07692};
        11'd  833 , 11'd 1327 : sin_data <= {-16'd07755};
        11'd  834 , 11'd 1326 : sin_data <= {-16'd07818};
        11'd  835 , 11'd 1325 : sin_data <= {-16'd07881};
        11'd  836 , 11'd 1324 : sin_data <= {-16'd07943};
        11'd  837 , 11'd 1323 : sin_data <= {-16'd08006};
        11'd  838 , 11'd 1322 : sin_data <= {-16'd08068};
        11'd  839 , 11'd 1321 : sin_data <= {-16'd08130};
        11'd  840 , 11'd 1320 : sin_data <= {-16'd08192};
        11'd  841 , 11'd 1319 : sin_data <= {-16'd08254};
        11'd  842 , 11'd 1318 : sin_data <= {-16'd08316};
        11'd  843 , 11'd 1317 : sin_data <= {-16'd08377};
        11'd  844 , 11'd 1316 : sin_data <= {-16'd08438};
        11'd  845 , 11'd 1315 : sin_data <= {-16'd08500};
        11'd  846 , 11'd 1314 : sin_data <= {-16'd08561};
        11'd  847 , 11'd 1313 : sin_data <= {-16'd08621};
        11'd  848 , 11'd 1312 : sin_data <= {-16'd08682};
        11'd  849 , 11'd 1311 : sin_data <= {-16'd08743};
        11'd  850 , 11'd 1310 : sin_data <= {-16'd08803};
        11'd  851 , 11'd 1309 : sin_data <= {-16'd08863};
        11'd  852 , 11'd 1308 : sin_data <= {-16'd08923};
        11'd  853 , 11'd 1307 : sin_data <= {-16'd08983};
        11'd  854 , 11'd 1306 : sin_data <= {-16'd09043};
        11'd  855 , 11'd 1305 : sin_data <= {-16'd09102};
        11'd  856 , 11'd 1304 : sin_data <= {-16'd09162};
        11'd  857 , 11'd 1303 : sin_data <= {-16'd09221};
        11'd  858 , 11'd 1302 : sin_data <= {-16'd09280};
        11'd  859 , 11'd 1301 : sin_data <= {-16'd09339};
        11'd  860 , 11'd 1300 : sin_data <= {-16'd09397};
        11'd  861 , 11'd 1299 : sin_data <= {-16'd09456};
        11'd  862 , 11'd 1298 : sin_data <= {-16'd09514};
        11'd  863 , 11'd 1297 : sin_data <= {-16'd09572};
        11'd  864 , 11'd 1296 : sin_data <= {-16'd09630};
        11'd  865 , 11'd 1295 : sin_data <= {-16'd09688};
        11'd  866 , 11'd 1294 : sin_data <= {-16'd09746};
        11'd  867 , 11'd 1293 : sin_data <= {-16'd09803};
        11'd  868 , 11'd 1292 : sin_data <= {-16'd09860};
        11'd  869 , 11'd 1291 : sin_data <= {-16'd09917};
        11'd  870 , 11'd 1290 : sin_data <= {-16'd09974};
        11'd  871 , 11'd 1289 : sin_data <= {-16'd10031};
        11'd  872 , 11'd 1288 : sin_data <= {-16'd10087};
        11'd  873 , 11'd 1287 : sin_data <= {-16'd10143};
        11'd  874 , 11'd 1286 : sin_data <= {-16'd10199};
        11'd  875 , 11'd 1285 : sin_data <= {-16'd10255};
        11'd  876 , 11'd 1284 : sin_data <= {-16'd10311};
        11'd  877 , 11'd 1283 : sin_data <= {-16'd10366};
        11'd  878 , 11'd 1282 : sin_data <= {-16'd10422};
        11'd  879 , 11'd 1281 : sin_data <= {-16'd10477};
        11'd  880 , 11'd 1280 : sin_data <= {-16'd10531};
        11'd  881 , 11'd 1279 : sin_data <= {-16'd10586};
        11'd  882 , 11'd 1278 : sin_data <= {-16'd10641};
        11'd  883 , 11'd 1277 : sin_data <= {-16'd10695};
        11'd  884 , 11'd 1276 : sin_data <= {-16'd10749};
        11'd  885 , 11'd 1275 : sin_data <= {-16'd10803};
        11'd  886 , 11'd 1274 : sin_data <= {-16'd10856};
        11'd  887 , 11'd 1273 : sin_data <= {-16'd10910};
        11'd  888 , 11'd 1272 : sin_data <= {-16'd10963};
        11'd  889 , 11'd 1271 : sin_data <= {-16'd11016};
        11'd  890 , 11'd 1270 : sin_data <= {-16'd11069};
        11'd  891 , 11'd 1269 : sin_data <= {-16'd11121};
        11'd  892 , 11'd 1268 : sin_data <= {-16'd11174};
        11'd  893 , 11'd 1267 : sin_data <= {-16'd11226};
        11'd  894 , 11'd 1266 : sin_data <= {-16'd11278};
        11'd  895 , 11'd 1265 : sin_data <= {-16'd11330};
        11'd  896 , 11'd 1264 : sin_data <= {-16'd11381};
        11'd  897 , 11'd 1263 : sin_data <= {-16'd11433};
        11'd  898 , 11'd 1262 : sin_data <= {-16'd11484};
        11'd  899 , 11'd 1261 : sin_data <= {-16'd11535};
        11'd  900 , 11'd 1260 : sin_data <= {-16'd11585};
        11'd  901 , 11'd 1259 : sin_data <= {-16'd11636};
        11'd  902 , 11'd 1258 : sin_data <= {-16'd11686};
        11'd  903 , 11'd 1257 : sin_data <= {-16'd11736};
        11'd  904 , 11'd 1256 : sin_data <= {-16'd11786};
        11'd  905 , 11'd 1255 : sin_data <= {-16'd11835};
        11'd  906 , 11'd 1254 : sin_data <= {-16'd11885};
        11'd  907 , 11'd 1253 : sin_data <= {-16'd11934};
        11'd  908 , 11'd 1252 : sin_data <= {-16'd11982};
        11'd  909 , 11'd 1251 : sin_data <= {-16'd12031};
        11'd  910 , 11'd 1250 : sin_data <= {-16'd12080};
        11'd  911 , 11'd 1249 : sin_data <= {-16'd12128};
        11'd  912 , 11'd 1248 : sin_data <= {-16'd12176};
        11'd  913 , 11'd 1247 : sin_data <= {-16'd12223};
        11'd  914 , 11'd 1246 : sin_data <= {-16'd12271};
        11'd  915 , 11'd 1245 : sin_data <= {-16'd12318};
        11'd  916 , 11'd 1244 : sin_data <= {-16'd12365};
        11'd  917 , 11'd 1243 : sin_data <= {-16'd12412};
        11'd  918 , 11'd 1242 : sin_data <= {-16'd12458};
        11'd  919 , 11'd 1241 : sin_data <= {-16'd12505};
        11'd  920 , 11'd 1240 : sin_data <= {-16'd12551};
        11'd  921 , 11'd 1239 : sin_data <= {-16'd12597};
        11'd  922 , 11'd 1238 : sin_data <= {-16'd12642};
        11'd  923 , 11'd 1237 : sin_data <= {-16'd12688};
        11'd  924 , 11'd 1236 : sin_data <= {-16'd12733};
        11'd  925 , 11'd 1235 : sin_data <= {-16'd12778};
        11'd  926 , 11'd 1234 : sin_data <= {-16'd12822};
        11'd  927 , 11'd 1233 : sin_data <= {-16'd12867};
        11'd  928 , 11'd 1232 : sin_data <= {-16'd12911};
        11'd  929 , 11'd 1231 : sin_data <= {-16'd12955};
        11'd  930 , 11'd 1230 : sin_data <= {-16'd12998};
        11'd  931 , 11'd 1229 : sin_data <= {-16'd13042};
        11'd  932 , 11'd 1228 : sin_data <= {-16'd13085};
        11'd  933 , 11'd 1227 : sin_data <= {-16'd13128};
        11'd  934 , 11'd 1226 : sin_data <= {-16'd13170};
        11'd  935 , 11'd 1225 : sin_data <= {-16'd13213};
        11'd  936 , 11'd 1224 : sin_data <= {-16'd13255};
        11'd  937 , 11'd 1223 : sin_data <= {-16'd13297};
        11'd  938 , 11'd 1222 : sin_data <= {-16'd13338};
        11'd  939 , 11'd 1221 : sin_data <= {-16'd13380};
        11'd  940 , 11'd 1220 : sin_data <= {-16'd13421};
        11'd  941 , 11'd 1219 : sin_data <= {-16'd13462};
        11'd  942 , 11'd 1218 : sin_data <= {-16'd13502};
        11'd  943 , 11'd 1217 : sin_data <= {-16'd13543};
        11'd  944 , 11'd 1216 : sin_data <= {-16'd13583};
        11'd  945 , 11'd 1215 : sin_data <= {-16'd13623};
        11'd  946 , 11'd 1214 : sin_data <= {-16'd13662};
        11'd  947 , 11'd 1213 : sin_data <= {-16'd13702};
        11'd  948 , 11'd 1212 : sin_data <= {-16'd13741};
        11'd  949 , 11'd 1211 : sin_data <= {-16'd13780};
        11'd  950 , 11'd 1210 : sin_data <= {-16'd13818};
        11'd  951 , 11'd 1209 : sin_data <= {-16'd13856};
        11'd  952 , 11'd 1208 : sin_data <= {-16'd13894};
        11'd  953 , 11'd 1207 : sin_data <= {-16'd13932};
        11'd  954 , 11'd 1206 : sin_data <= {-16'd13970};
        11'd  955 , 11'd 1205 : sin_data <= {-16'd14007};
        11'd  956 , 11'd 1204 : sin_data <= {-16'd14044};
        11'd  957 , 11'd 1203 : sin_data <= {-16'd14081};
        11'd  958 , 11'd 1202 : sin_data <= {-16'd14117};
        11'd  959 , 11'd 1201 : sin_data <= {-16'd14153};
        11'd  960 , 11'd 1200 : sin_data <= {-16'd14189};
        11'd  961 , 11'd 1199 : sin_data <= {-16'd14225};
        11'd  962 , 11'd 1198 : sin_data <= {-16'd14260};
        11'd  963 , 11'd 1197 : sin_data <= {-16'd14295};
        11'd  964 , 11'd 1196 : sin_data <= {-16'd14330};
        11'd  965 , 11'd 1195 : sin_data <= {-16'd14364};
        11'd  966 , 11'd 1194 : sin_data <= {-16'd14399};
        11'd  967 , 11'd 1193 : sin_data <= {-16'd14433};
        11'd  968 , 11'd 1192 : sin_data <= {-16'd14466};
        11'd  969 , 11'd 1191 : sin_data <= {-16'd14500};
        11'd  970 , 11'd 1190 : sin_data <= {-16'd14533};
        11'd  971 , 11'd 1189 : sin_data <= {-16'd14566};
        11'd  972 , 11'd 1188 : sin_data <= {-16'd14598};
        11'd  973 , 11'd 1187 : sin_data <= {-16'd14631};
        11'd  974 , 11'd 1186 : sin_data <= {-16'd14663};
        11'd  975 , 11'd 1185 : sin_data <= {-16'd14694};
        11'd  976 , 11'd 1184 : sin_data <= {-16'd14726};
        11'd  977 , 11'd 1183 : sin_data <= {-16'd14757};
        11'd  978 , 11'd 1182 : sin_data <= {-16'd14788};
        11'd  979 , 11'd 1181 : sin_data <= {-16'd14819};
        11'd  980 , 11'd 1180 : sin_data <= {-16'd14849};
        11'd  981 , 11'd 1179 : sin_data <= {-16'd14879};
        11'd  982 , 11'd 1178 : sin_data <= {-16'd14909};
        11'd  983 , 11'd 1177 : sin_data <= {-16'd14938};
        11'd  984 , 11'd 1176 : sin_data <= {-16'd14968};
        11'd  985 , 11'd 1175 : sin_data <= {-16'd14996};
        11'd  986 , 11'd 1174 : sin_data <= {-16'd15025};
        11'd  987 , 11'd 1173 : sin_data <= {-16'd15053};
        11'd  988 , 11'd 1172 : sin_data <= {-16'd15082};
        11'd  989 , 11'd 1171 : sin_data <= {-16'd15109};
        11'd  990 , 11'd 1170 : sin_data <= {-16'd15137};
        11'd  991 , 11'd 1169 : sin_data <= {-16'd15164};
        11'd  992 , 11'd 1168 : sin_data <= {-16'd15191};
        11'd  993 , 11'd 1167 : sin_data <= {-16'd15218};
        11'd  994 , 11'd 1166 : sin_data <= {-16'd15244};
        11'd  995 , 11'd 1165 : sin_data <= {-16'd15270};
        11'd  996 , 11'd 1164 : sin_data <= {-16'd15296};
        11'd  997 , 11'd 1163 : sin_data <= {-16'd15321};
        11'd  998 , 11'd 1162 : sin_data <= {-16'd15346};
        11'd  999 , 11'd 1161 : sin_data <= {-16'd15371};
        11'd 1000 , 11'd 1160 : sin_data <= {-16'd15396};
        11'd 1001 , 11'd 1159 : sin_data <= {-16'd15420};
        11'd 1002 , 11'd 1158 : sin_data <= {-16'd15444};
        11'd 1003 , 11'd 1157 : sin_data <= {-16'd15468};
        11'd 1004 , 11'd 1156 : sin_data <= {-16'd15491};
        11'd 1005 , 11'd 1155 : sin_data <= {-16'd15515};
        11'd 1006 , 11'd 1154 : sin_data <= {-16'd15537};
        11'd 1007 , 11'd 1153 : sin_data <= {-16'd15560};
        11'd 1008 , 11'd 1152 : sin_data <= {-16'd15582};
        11'd 1009 , 11'd 1151 : sin_data <= {-16'd15604};
        11'd 1010 , 11'd 1150 : sin_data <= {-16'd15626};
        11'd 1011 , 11'd 1149 : sin_data <= {-16'd15647};
        11'd 1012 , 11'd 1148 : sin_data <= {-16'd15668};
        11'd 1013 , 11'd 1147 : sin_data <= {-16'd15689};
        11'd 1014 , 11'd 1146 : sin_data <= {-16'd15709};
        11'd 1015 , 11'd 1145 : sin_data <= {-16'd15729};
        11'd 1016 , 11'd 1144 : sin_data <= {-16'd15749};
        11'd 1017 , 11'd 1143 : sin_data <= {-16'd15769};
        11'd 1018 , 11'd 1142 : sin_data <= {-16'd15788};
        11'd 1019 , 11'd 1141 : sin_data <= {-16'd15807};
        11'd 1020 , 11'd 1140 : sin_data <= {-16'd15826};
        11'd 1021 , 11'd 1139 : sin_data <= {-16'd15844};
        11'd 1022 , 11'd 1138 : sin_data <= {-16'd15862};
        11'd 1023 , 11'd 1137 : sin_data <= {-16'd15880};
        11'd 1024 , 11'd 1136 : sin_data <= {-16'd15897};
        11'd 1025 , 11'd 1135 : sin_data <= {-16'd15914};
        11'd 1026 , 11'd 1134 : sin_data <= {-16'd15931};
        11'd 1027 , 11'd 1133 : sin_data <= {-16'd15948};
        11'd 1028 , 11'd 1132 : sin_data <= {-16'd15964};
        11'd 1029 , 11'd 1131 : sin_data <= {-16'd15980};
        11'd 1030 , 11'd 1130 : sin_data <= {-16'd15996};
        11'd 1031 , 11'd 1129 : sin_data <= {-16'd16011};
        11'd 1032 , 11'd 1128 : sin_data <= {-16'd16026};
        11'd 1033 , 11'd 1127 : sin_data <= {-16'd16041};
        11'd 1034 , 11'd 1126 : sin_data <= {-16'd16055};
        11'd 1035 , 11'd 1125 : sin_data <= {-16'd16069};
        11'd 1036 , 11'd 1124 : sin_data <= {-16'd16083};
        11'd 1037 , 11'd 1123 : sin_data <= {-16'd16096};
        11'd 1038 , 11'd 1122 : sin_data <= {-16'd16110};
        11'd 1039 , 11'd 1121 : sin_data <= {-16'd16123};
        11'd 1040 , 11'd 1120 : sin_data <= {-16'd16135};
        11'd 1041 , 11'd 1119 : sin_data <= {-16'd16147};
        11'd 1042 , 11'd 1118 : sin_data <= {-16'd16159};
        11'd 1043 , 11'd 1117 : sin_data <= {-16'd16171};
        11'd 1044 , 11'd 1116 : sin_data <= {-16'd16182};
        11'd 1045 , 11'd 1115 : sin_data <= {-16'd16193};
        11'd 1046 , 11'd 1114 : sin_data <= {-16'd16204};
        11'd 1047 , 11'd 1113 : sin_data <= {-16'd16214};
        11'd 1048 , 11'd 1112 : sin_data <= {-16'd16225};
        11'd 1049 , 11'd 1111 : sin_data <= {-16'd16234};
        11'd 1050 , 11'd 1110 : sin_data <= {-16'd16244};
        11'd 1051 , 11'd 1109 : sin_data <= {-16'd16253};
        11'd 1052 , 11'd 1108 : sin_data <= {-16'd16262};
        11'd 1053 , 11'd 1107 : sin_data <= {-16'd16270};
        11'd 1054 , 11'd 1106 : sin_data <= {-16'd16279};
        11'd 1055 , 11'd 1105 : sin_data <= {-16'd16287};
        11'd 1056 , 11'd 1104 : sin_data <= {-16'd16294};
        11'd 1057 , 11'd 1103 : sin_data <= {-16'd16302};
        11'd 1058 , 11'd 1102 : sin_data <= {-16'd16309};
        11'd 1059 , 11'd 1101 : sin_data <= {-16'd16315};
        11'd 1060 , 11'd 1100 : sin_data <= {-16'd16322};
        11'd 1061 , 11'd 1099 : sin_data <= {-16'd16328};
        11'd 1062 , 11'd 1098 : sin_data <= {-16'd16333};
        11'd 1063 , 11'd 1097 : sin_data <= {-16'd16339};
        11'd 1064 , 11'd 1096 : sin_data <= {-16'd16344};
        11'd 1065 , 11'd 1095 : sin_data <= {-16'd16349};
        11'd 1066 , 11'd 1094 : sin_data <= {-16'd16353};
        11'd 1067 , 11'd 1093 : sin_data <= {-16'd16358};
        11'd 1068 , 11'd 1092 : sin_data <= {-16'd16362};
        11'd 1069 , 11'd 1091 : sin_data <= {-16'd16365};
        11'd 1070 , 11'd 1090 : sin_data <= {-16'd16368};
        11'd 1071 , 11'd 1089 : sin_data <= {-16'd16371};
        11'd 1072 , 11'd 1088 : sin_data <= {-16'd16374};
        11'd 1073 , 11'd 1087 : sin_data <= {-16'd16376};
        11'd 1074 , 11'd 1086 : sin_data <= {-16'd16378};
        11'd 1075 , 11'd 1085 : sin_data <= {-16'd16380};
        11'd 1076 , 11'd 1084 : sin_data <= {-16'd16382};
        11'd 1077 , 11'd 1083 : sin_data <= {-16'd16383};
        11'd 1078 , 11'd 1082 : sin_data <= {-16'd16383};
        11'd 1079 , 11'd 1081 : sin_data <= {-16'd16384};
        11'd 1080             : sin_data <= {-16'd16384};
        
        default: sin_data <= {16'd0000};
    endcase
end

always@(angle_div4) begin
    case(angle_div4)
        11'd    0 , 11'd 1440 : cos_data <= {16'd16384};
        11'd    1 , 11'd 1439 : cos_data <= {16'd16384};
        11'd    2 , 11'd 1438 : cos_data <= {16'd16383};
        11'd    3 , 11'd 1437 : cos_data <= {16'd16383};
        11'd    4 , 11'd 1436 : cos_data <= {16'd16382};
        11'd    5 , 11'd 1435 : cos_data <= {16'd16380};
        11'd    6 , 11'd 1434 : cos_data <= {16'd16378};
        11'd    7 , 11'd 1433 : cos_data <= {16'd16376};
        11'd    8 , 11'd 1432 : cos_data <= {16'd16374};
        11'd    9 , 11'd 1431 : cos_data <= {16'd16371};
        11'd   10 , 11'd 1430 : cos_data <= {16'd16368};
        11'd   11 , 11'd 1429 : cos_data <= {16'd16365};
        11'd   12 , 11'd 1428 : cos_data <= {16'd16362};
        11'd   13 , 11'd 1427 : cos_data <= {16'd16358};
        11'd   14 , 11'd 1426 : cos_data <= {16'd16353};
        11'd   15 , 11'd 1425 : cos_data <= {16'd16349};
        11'd   16 , 11'd 1424 : cos_data <= {16'd16344};
        11'd   17 , 11'd 1423 : cos_data <= {16'd16339};
        11'd   18 , 11'd 1422 : cos_data <= {16'd16333};
        11'd   19 , 11'd 1421 : cos_data <= {16'd16328};
        11'd   20 , 11'd 1420 : cos_data <= {16'd16322};
        11'd   21 , 11'd 1419 : cos_data <= {16'd16315};
        11'd   22 , 11'd 1418 : cos_data <= {16'd16309};
        11'd   23 , 11'd 1417 : cos_data <= {16'd16302};
        11'd   24 , 11'd 1416 : cos_data <= {16'd16294};
        11'd   25 , 11'd 1415 : cos_data <= {16'd16287};
        11'd   26 , 11'd 1414 : cos_data <= {16'd16279};
        11'd   27 , 11'd 1413 : cos_data <= {16'd16270};
        11'd   28 , 11'd 1412 : cos_data <= {16'd16262};
        11'd   29 , 11'd 1411 : cos_data <= {16'd16253};
        11'd   30 , 11'd 1410 : cos_data <= {16'd16244};
        11'd   31 , 11'd 1409 : cos_data <= {16'd16234};
        11'd   32 , 11'd 1408 : cos_data <= {16'd16225};
        11'd   33 , 11'd 1407 : cos_data <= {16'd16214};
        11'd   34 , 11'd 1406 : cos_data <= {16'd16204};
        11'd   35 , 11'd 1405 : cos_data <= {16'd16193};
        11'd   36 , 11'd 1404 : cos_data <= {16'd16182};
        11'd   37 , 11'd 1403 : cos_data <= {16'd16171};
        11'd   38 , 11'd 1402 : cos_data <= {16'd16159};
        11'd   39 , 11'd 1401 : cos_data <= {16'd16147};
        11'd   40 , 11'd 1400 : cos_data <= {16'd16135};
        11'd   41 , 11'd 1399 : cos_data <= {16'd16123};
        11'd   42 , 11'd 1398 : cos_data <= {16'd16110};
        11'd   43 , 11'd 1397 : cos_data <= {16'd16096};
        11'd   44 , 11'd 1396 : cos_data <= {16'd16083};
        11'd   45 , 11'd 1395 : cos_data <= {16'd16069};
        11'd   46 , 11'd 1394 : cos_data <= {16'd16055};
        11'd   47 , 11'd 1393 : cos_data <= {16'd16041};
        11'd   48 , 11'd 1392 : cos_data <= {16'd16026};
        11'd   49 , 11'd 1391 : cos_data <= {16'd16011};
        11'd   50 , 11'd 1390 : cos_data <= {16'd15996};
        11'd   51 , 11'd 1389 : cos_data <= {16'd15980};
        11'd   52 , 11'd 1388 : cos_data <= {16'd15964};
        11'd   53 , 11'd 1387 : cos_data <= {16'd15948};
        11'd   54 , 11'd 1386 : cos_data <= {16'd15931};
        11'd   55 , 11'd 1385 : cos_data <= {16'd15914};
        11'd   56 , 11'd 1384 : cos_data <= {16'd15897};
        11'd   57 , 11'd 1383 : cos_data <= {16'd15880};
        11'd   58 , 11'd 1382 : cos_data <= {16'd15862};
        11'd   59 , 11'd 1381 : cos_data <= {16'd15844};
        11'd   60 , 11'd 1380 : cos_data <= {16'd15826};
        11'd   61 , 11'd 1379 : cos_data <= {16'd15807};
        11'd   62 , 11'd 1378 : cos_data <= {16'd15788};
        11'd   63 , 11'd 1377 : cos_data <= {16'd15769};
        11'd   64 , 11'd 1376 : cos_data <= {16'd15749};
        11'd   65 , 11'd 1375 : cos_data <= {16'd15729};
        11'd   66 , 11'd 1374 : cos_data <= {16'd15709};
        11'd   67 , 11'd 1373 : cos_data <= {16'd15689};
        11'd   68 , 11'd 1372 : cos_data <= {16'd15668};
        11'd   69 , 11'd 1371 : cos_data <= {16'd15647};
        11'd   70 , 11'd 1370 : cos_data <= {16'd15626};
        11'd   71 , 11'd 1369 : cos_data <= {16'd15604};
        11'd   72 , 11'd 1368 : cos_data <= {16'd15582};
        11'd   73 , 11'd 1367 : cos_data <= {16'd15560};
        11'd   74 , 11'd 1366 : cos_data <= {16'd15537};
        11'd   75 , 11'd 1365 : cos_data <= {16'd15515};
        11'd   76 , 11'd 1364 : cos_data <= {16'd15491};
        11'd   77 , 11'd 1363 : cos_data <= {16'd15468};
        11'd   78 , 11'd 1362 : cos_data <= {16'd15444};
        11'd   79 , 11'd 1361 : cos_data <= {16'd15420};
        11'd   80 , 11'd 1360 : cos_data <= {16'd15396};
        11'd   81 , 11'd 1359 : cos_data <= {16'd15371};
        11'd   82 , 11'd 1358 : cos_data <= {16'd15346};
        11'd   83 , 11'd 1357 : cos_data <= {16'd15321};
        11'd   84 , 11'd 1356 : cos_data <= {16'd15296};
        11'd   85 , 11'd 1355 : cos_data <= {16'd15270};
        11'd   86 , 11'd 1354 : cos_data <= {16'd15244};
        11'd   87 , 11'd 1353 : cos_data <= {16'd15218};
        11'd   88 , 11'd 1352 : cos_data <= {16'd15191};
        11'd   89 , 11'd 1351 : cos_data <= {16'd15164};
        11'd   90 , 11'd 1350 : cos_data <= {16'd15137};
        11'd   91 , 11'd 1349 : cos_data <= {16'd15109};
        11'd   92 , 11'd 1348 : cos_data <= {16'd15082};
        11'd   93 , 11'd 1347 : cos_data <= {16'd15053};
        11'd   94 , 11'd 1346 : cos_data <= {16'd15025};
        11'd   95 , 11'd 1345 : cos_data <= {16'd14996};
        11'd   96 , 11'd 1344 : cos_data <= {16'd14968};
        11'd   97 , 11'd 1343 : cos_data <= {16'd14938};
        11'd   98 , 11'd 1342 : cos_data <= {16'd14909};
        11'd   99 , 11'd 1341 : cos_data <= {16'd14879};
        11'd  100 , 11'd 1340 : cos_data <= {16'd14849};
        11'd  101 , 11'd 1339 : cos_data <= {16'd14819};
        11'd  102 , 11'd 1338 : cos_data <= {16'd14788};
        11'd  103 , 11'd 1337 : cos_data <= {16'd14757};
        11'd  104 , 11'd 1336 : cos_data <= {16'd14726};
        11'd  105 , 11'd 1335 : cos_data <= {16'd14694};
        11'd  106 , 11'd 1334 : cos_data <= {16'd14663};
        11'd  107 , 11'd 1333 : cos_data <= {16'd14631};
        11'd  108 , 11'd 1332 : cos_data <= {16'd14598};
        11'd  109 , 11'd 1331 : cos_data <= {16'd14566};
        11'd  110 , 11'd 1330 : cos_data <= {16'd14533};
        11'd  111 , 11'd 1329 : cos_data <= {16'd14500};
        11'd  112 , 11'd 1328 : cos_data <= {16'd14466};
        11'd  113 , 11'd 1327 : cos_data <= {16'd14433};
        11'd  114 , 11'd 1326 : cos_data <= {16'd14399};
        11'd  115 , 11'd 1325 : cos_data <= {16'd14364};
        11'd  116 , 11'd 1324 : cos_data <= {16'd14330};
        11'd  117 , 11'd 1323 : cos_data <= {16'd14295};
        11'd  118 , 11'd 1322 : cos_data <= {16'd14260};
        11'd  119 , 11'd 1321 : cos_data <= {16'd14225};
        11'd  120 , 11'd 1320 : cos_data <= {16'd14189};
        11'd  121 , 11'd 1319 : cos_data <= {16'd14153};
        11'd  122 , 11'd 1318 : cos_data <= {16'd14117};
        11'd  123 , 11'd 1317 : cos_data <= {16'd14081};
        11'd  124 , 11'd 1316 : cos_data <= {16'd14044};
        11'd  125 , 11'd 1315 : cos_data <= {16'd14007};
        11'd  126 , 11'd 1314 : cos_data <= {16'd13970};
        11'd  127 , 11'd 1313 : cos_data <= {16'd13932};
        11'd  128 , 11'd 1312 : cos_data <= {16'd13894};
        11'd  129 , 11'd 1311 : cos_data <= {16'd13856};
        11'd  130 , 11'd 1310 : cos_data <= {16'd13818};
        11'd  131 , 11'd 1309 : cos_data <= {16'd13780};
        11'd  132 , 11'd 1308 : cos_data <= {16'd13741};
        11'd  133 , 11'd 1307 : cos_data <= {16'd13702};
        11'd  134 , 11'd 1306 : cos_data <= {16'd13662};
        11'd  135 , 11'd 1305 : cos_data <= {16'd13623};
        11'd  136 , 11'd 1304 : cos_data <= {16'd13583};
        11'd  137 , 11'd 1303 : cos_data <= {16'd13543};
        11'd  138 , 11'd 1302 : cos_data <= {16'd13502};
        11'd  139 , 11'd 1301 : cos_data <= {16'd13462};
        11'd  140 , 11'd 1300 : cos_data <= {16'd13421};
        11'd  141 , 11'd 1299 : cos_data <= {16'd13380};
        11'd  142 , 11'd 1298 : cos_data <= {16'd13338};
        11'd  143 , 11'd 1297 : cos_data <= {16'd13297};
        11'd  144 , 11'd 1296 : cos_data <= {16'd13255};
        11'd  145 , 11'd 1295 : cos_data <= {16'd13213};
        11'd  146 , 11'd 1294 : cos_data <= {16'd13170};
        11'd  147 , 11'd 1293 : cos_data <= {16'd13128};
        11'd  148 , 11'd 1292 : cos_data <= {16'd13085};
        11'd  149 , 11'd 1291 : cos_data <= {16'd13042};
        11'd  150 , 11'd 1290 : cos_data <= {16'd12998};
        11'd  151 , 11'd 1289 : cos_data <= {16'd12955};
        11'd  152 , 11'd 1288 : cos_data <= {16'd12911};
        11'd  153 , 11'd 1287 : cos_data <= {16'd12867};
        11'd  154 , 11'd 1286 : cos_data <= {16'd12822};
        11'd  155 , 11'd 1285 : cos_data <= {16'd12778};
        11'd  156 , 11'd 1284 : cos_data <= {16'd12733};
        11'd  157 , 11'd 1283 : cos_data <= {16'd12688};
        11'd  158 , 11'd 1282 : cos_data <= {16'd12642};
        11'd  159 , 11'd 1281 : cos_data <= {16'd12597};
        11'd  160 , 11'd 1280 : cos_data <= {16'd12551};
        11'd  161 , 11'd 1279 : cos_data <= {16'd12505};
        11'd  162 , 11'd 1278 : cos_data <= {16'd12458};
        11'd  163 , 11'd 1277 : cos_data <= {16'd12412};
        11'd  164 , 11'd 1276 : cos_data <= {16'd12365};
        11'd  165 , 11'd 1275 : cos_data <= {16'd12318};
        11'd  166 , 11'd 1274 : cos_data <= {16'd12271};
        11'd  167 , 11'd 1273 : cos_data <= {16'd12223};
        11'd  168 , 11'd 1272 : cos_data <= {16'd12176};
        11'd  169 , 11'd 1271 : cos_data <= {16'd12128};
        11'd  170 , 11'd 1270 : cos_data <= {16'd12080};
        11'd  171 , 11'd 1269 : cos_data <= {16'd12031};
        11'd  172 , 11'd 1268 : cos_data <= {16'd11982};
        11'd  173 , 11'd 1267 : cos_data <= {16'd11934};
        11'd  174 , 11'd 1266 : cos_data <= {16'd11885};
        11'd  175 , 11'd 1265 : cos_data <= {16'd11835};
        11'd  176 , 11'd 1264 : cos_data <= {16'd11786};
        11'd  177 , 11'd 1263 : cos_data <= {16'd11736};
        11'd  178 , 11'd 1262 : cos_data <= {16'd11686};
        11'd  179 , 11'd 1261 : cos_data <= {16'd11636};
        11'd  180 , 11'd 1260 : cos_data <= {16'd11585};
        11'd  181 , 11'd 1259 : cos_data <= {16'd11535};
        11'd  182 , 11'd 1258 : cos_data <= {16'd11484};
        11'd  183 , 11'd 1257 : cos_data <= {16'd11433};
        11'd  184 , 11'd 1256 : cos_data <= {16'd11381};
        11'd  185 , 11'd 1255 : cos_data <= {16'd11330};
        11'd  186 , 11'd 1254 : cos_data <= {16'd11278};
        11'd  187 , 11'd 1253 : cos_data <= {16'd11226};
        11'd  188 , 11'd 1252 : cos_data <= {16'd11174};
        11'd  189 , 11'd 1251 : cos_data <= {16'd11121};
        11'd  190 , 11'd 1250 : cos_data <= {16'd11069};
        11'd  191 , 11'd 1249 : cos_data <= {16'd11016};
        11'd  192 , 11'd 1248 : cos_data <= {16'd10963};
        11'd  193 , 11'd 1247 : cos_data <= {16'd10910};
        11'd  194 , 11'd 1246 : cos_data <= {16'd10856};
        11'd  195 , 11'd 1245 : cos_data <= {16'd10803};
        11'd  196 , 11'd 1244 : cos_data <= {16'd10749};
        11'd  197 , 11'd 1243 : cos_data <= {16'd10695};
        11'd  198 , 11'd 1242 : cos_data <= {16'd10641};
        11'd  199 , 11'd 1241 : cos_data <= {16'd10586};
        11'd  200 , 11'd 1240 : cos_data <= {16'd10531};
        11'd  201 , 11'd 1239 : cos_data <= {16'd10477};
        11'd  202 , 11'd 1238 : cos_data <= {16'd10422};
        11'd  203 , 11'd 1237 : cos_data <= {16'd10366};
        11'd  204 , 11'd 1236 : cos_data <= {16'd10311};
        11'd  205 , 11'd 1235 : cos_data <= {16'd10255};
        11'd  206 , 11'd 1234 : cos_data <= {16'd10199};
        11'd  207 , 11'd 1233 : cos_data <= {16'd10143};
        11'd  208 , 11'd 1232 : cos_data <= {16'd10087};
        11'd  209 , 11'd 1231 : cos_data <= {16'd10031};
        11'd  210 , 11'd 1230 : cos_data <= {16'd09974};
        11'd  211 , 11'd 1229 : cos_data <= {16'd09917};
        11'd  212 , 11'd 1228 : cos_data <= {16'd09860};
        11'd  213 , 11'd 1227 : cos_data <= {16'd09803};
        11'd  214 , 11'd 1226 : cos_data <= {16'd09746};
        11'd  215 , 11'd 1225 : cos_data <= {16'd09688};
        11'd  216 , 11'd 1224 : cos_data <= {16'd09630};
        11'd  217 , 11'd 1223 : cos_data <= {16'd09572};
        11'd  218 , 11'd 1222 : cos_data <= {16'd09514};
        11'd  219 , 11'd 1221 : cos_data <= {16'd09456};
        11'd  220 , 11'd 1220 : cos_data <= {16'd09397};
        11'd  221 , 11'd 1219 : cos_data <= {16'd09339};
        11'd  222 , 11'd 1218 : cos_data <= {16'd09280};
        11'd  223 , 11'd 1217 : cos_data <= {16'd09221};
        11'd  224 , 11'd 1216 : cos_data <= {16'd09162};
        11'd  225 , 11'd 1215 : cos_data <= {16'd09102};
        11'd  226 , 11'd 1214 : cos_data <= {16'd09043};
        11'd  227 , 11'd 1213 : cos_data <= {16'd08983};
        11'd  228 , 11'd 1212 : cos_data <= {16'd08923};
        11'd  229 , 11'd 1211 : cos_data <= {16'd08863};
        11'd  230 , 11'd 1210 : cos_data <= {16'd08803};
        11'd  231 , 11'd 1209 : cos_data <= {16'd08743};
        11'd  232 , 11'd 1208 : cos_data <= {16'd08682};
        11'd  233 , 11'd 1207 : cos_data <= {16'd08621};
        11'd  234 , 11'd 1206 : cos_data <= {16'd08561};
        11'd  235 , 11'd 1205 : cos_data <= {16'd08500};
        11'd  236 , 11'd 1204 : cos_data <= {16'd08438};
        11'd  237 , 11'd 1203 : cos_data <= {16'd08377};
        11'd  238 , 11'd 1202 : cos_data <= {16'd08316};
        11'd  239 , 11'd 1201 : cos_data <= {16'd08254};
        11'd  240 , 11'd 1200 : cos_data <= {16'd08192};
        11'd  241 , 11'd 1199 : cos_data <= {16'd08130};
        11'd  242 , 11'd 1198 : cos_data <= {16'd08068};
        11'd  243 , 11'd 1197 : cos_data <= {16'd08006};
        11'd  244 , 11'd 1196 : cos_data <= {16'd07943};
        11'd  245 , 11'd 1195 : cos_data <= {16'd07881};
        11'd  246 , 11'd 1194 : cos_data <= {16'd07818};
        11'd  247 , 11'd 1193 : cos_data <= {16'd07755};
        11'd  248 , 11'd 1192 : cos_data <= {16'd07692};
        11'd  249 , 11'd 1191 : cos_data <= {16'd07629};
        11'd  250 , 11'd 1190 : cos_data <= {16'd07565};
        11'd  251 , 11'd 1189 : cos_data <= {16'd07502};
        11'd  252 , 11'd 1188 : cos_data <= {16'd07438};
        11'd  253 , 11'd 1187 : cos_data <= {16'd07374};
        11'd  254 , 11'd 1186 : cos_data <= {16'd07311};
        11'd  255 , 11'd 1185 : cos_data <= {16'd07246};
        11'd  256 , 11'd 1184 : cos_data <= {16'd07182};
        11'd  257 , 11'd 1183 : cos_data <= {16'd07118};
        11'd  258 , 11'd 1182 : cos_data <= {16'd07053};
        11'd  259 , 11'd 1181 : cos_data <= {16'd06989};
        11'd  260 , 11'd 1180 : cos_data <= {16'd06924};
        11'd  261 , 11'd 1179 : cos_data <= {16'd06859};
        11'd  262 , 11'd 1178 : cos_data <= {16'd06794};
        11'd  263 , 11'd 1177 : cos_data <= {16'd06729};
        11'd  264 , 11'd 1176 : cos_data <= {16'd06664};
        11'd  265 , 11'd 1175 : cos_data <= {16'd06599};
        11'd  266 , 11'd 1174 : cos_data <= {16'd06533};
        11'd  267 , 11'd 1173 : cos_data <= {16'd06467};
        11'd  268 , 11'd 1172 : cos_data <= {16'd06402};
        11'd  269 , 11'd 1171 : cos_data <= {16'd06336};
        11'd  270 , 11'd 1170 : cos_data <= {16'd06270};
        11'd  271 , 11'd 1169 : cos_data <= {16'd06204};
        11'd  272 , 11'd 1168 : cos_data <= {16'd06138};
        11'd  273 , 11'd 1167 : cos_data <= {16'd06071};
        11'd  274 , 11'd 1166 : cos_data <= {16'd06005};
        11'd  275 , 11'd 1165 : cos_data <= {16'd05938};
        11'd  276 , 11'd 1164 : cos_data <= {16'd05872};
        11'd  277 , 11'd 1163 : cos_data <= {16'd05805};
        11'd  278 , 11'd 1162 : cos_data <= {16'd05738};
        11'd  279 , 11'd 1161 : cos_data <= {16'd05671};
        11'd  280 , 11'd 1160 : cos_data <= {16'd05604};
        11'd  281 , 11'd 1159 : cos_data <= {16'd05536};
        11'd  282 , 11'd 1158 : cos_data <= {16'd05469};
        11'd  283 , 11'd 1157 : cos_data <= {16'd05402};
        11'd  284 , 11'd 1156 : cos_data <= {16'd05334};
        11'd  285 , 11'd 1155 : cos_data <= {16'd05266};
        11'd  286 , 11'd 1154 : cos_data <= {16'd05199};
        11'd  287 , 11'd 1153 : cos_data <= {16'd05131};
        11'd  288 , 11'd 1152 : cos_data <= {16'd05063};
        11'd  289 , 11'd 1151 : cos_data <= {16'd04995};
        11'd  290 , 11'd 1150 : cos_data <= {16'd04927};
        11'd  291 , 11'd 1149 : cos_data <= {16'd04859};
        11'd  292 , 11'd 1148 : cos_data <= {16'd04790};
        11'd  293 , 11'd 1147 : cos_data <= {16'd04722};
        11'd  294 , 11'd 1146 : cos_data <= {16'd04653};
        11'd  295 , 11'd 1145 : cos_data <= {16'd04585};
        11'd  296 , 11'd 1144 : cos_data <= {16'd04516};
        11'd  297 , 11'd 1143 : cos_data <= {16'd04447};
        11'd  298 , 11'd 1142 : cos_data <= {16'd04378};
        11'd  299 , 11'd 1141 : cos_data <= {16'd04310};
        11'd  300 , 11'd 1140 : cos_data <= {16'd04240};
        11'd  301 , 11'd 1139 : cos_data <= {16'd04171};
        11'd  302 , 11'd 1138 : cos_data <= {16'd04102};
        11'd  303 , 11'd 1137 : cos_data <= {16'd04033};
        11'd  304 , 11'd 1136 : cos_data <= {16'd03964};
        11'd  305 , 11'd 1135 : cos_data <= {16'd03894};
        11'd  306 , 11'd 1134 : cos_data <= {16'd03825};
        11'd  307 , 11'd 1133 : cos_data <= {16'd03755};
        11'd  308 , 11'd 1132 : cos_data <= {16'd03686};
        11'd  309 , 11'd 1131 : cos_data <= {16'd03616};
        11'd  310 , 11'd 1130 : cos_data <= {16'd03546};
        11'd  311 , 11'd 1129 : cos_data <= {16'd03476};
        11'd  312 , 11'd 1128 : cos_data <= {16'd03406};
        11'd  313 , 11'd 1127 : cos_data <= {16'd03336};
        11'd  314 , 11'd 1126 : cos_data <= {16'd03266};
        11'd  315 , 11'd 1125 : cos_data <= {16'd03196};
        11'd  316 , 11'd 1124 : cos_data <= {16'd03126};
        11'd  317 , 11'd 1123 : cos_data <= {16'd03056};
        11'd  318 , 11'd 1122 : cos_data <= {16'd02986};
        11'd  319 , 11'd 1121 : cos_data <= {16'd02915};
        11'd  320 , 11'd 1120 : cos_data <= {16'd02845};
        11'd  321 , 11'd 1119 : cos_data <= {16'd02775};
        11'd  322 , 11'd 1118 : cos_data <= {16'd02704};
        11'd  323 , 11'd 1117 : cos_data <= {16'd02634};
        11'd  324 , 11'd 1116 : cos_data <= {16'd02563};
        11'd  325 , 11'd 1115 : cos_data <= {16'd02492};
        11'd  326 , 11'd 1114 : cos_data <= {16'd02422};
        11'd  327 , 11'd 1113 : cos_data <= {16'd02351};
        11'd  328 , 11'd 1112 : cos_data <= {16'd02280};
        11'd  329 , 11'd 1111 : cos_data <= {16'd02209};
        11'd  330 , 11'd 1110 : cos_data <= {16'd02139};
        11'd  331 , 11'd 1109 : cos_data <= {16'd02068};
        11'd  332 , 11'd 1108 : cos_data <= {16'd01997};
        11'd  333 , 11'd 1107 : cos_data <= {16'd01926};
        11'd  334 , 11'd 1106 : cos_data <= {16'd01855};
        11'd  335 , 11'd 1105 : cos_data <= {16'd01784};
        11'd  336 , 11'd 1104 : cos_data <= {16'd01713};
        11'd  337 , 11'd 1103 : cos_data <= {16'd01641};
        11'd  338 , 11'd 1102 : cos_data <= {16'd01570};
        11'd  339 , 11'd 1101 : cos_data <= {16'd01499};
        11'd  340 , 11'd 1100 : cos_data <= {16'd01428};
        11'd  341 , 11'd 1099 : cos_data <= {16'd01357};
        11'd  342 , 11'd 1098 : cos_data <= {16'd01285};
        11'd  343 , 11'd 1097 : cos_data <= {16'd01214};
        11'd  344 , 11'd 1096 : cos_data <= {16'd01143};
        11'd  345 , 11'd 1095 : cos_data <= {16'd01072};
        11'd  346 , 11'd 1094 : cos_data <= {16'd01000};
        11'd  347 , 11'd 1093 : cos_data <= {16'd00929};
        11'd  348 , 11'd 1092 : cos_data <= {16'd00857};
        11'd  349 , 11'd 1091 : cos_data <= {16'd00786};
        11'd  350 , 11'd 1090 : cos_data <= {16'd00715};
        11'd  351 , 11'd 1089 : cos_data <= {16'd00643};
        11'd  352 , 11'd 1088 : cos_data <= {16'd00572};
        11'd  353 , 11'd 1087 : cos_data <= {16'd00500};
        11'd  354 , 11'd 1086 : cos_data <= {16'd00429};
        11'd  355 , 11'd 1085 : cos_data <= {16'd00357};
        11'd  356 , 11'd 1084 : cos_data <= {16'd00286};
        11'd  357 , 11'd 1083 : cos_data <= {16'd00214};
        11'd  358 , 11'd 1082 : cos_data <= {16'd00143};
        11'd  359 , 11'd 1081 : cos_data <= {16'd00071};
        11'd  360             : cos_data <= {16'd00000};
        



                   11'd 1080 : cos_data <= {-16'd00000};    
        11'd 361 , 11'd 1079 : cos_data <= {-16'd00071};
        11'd 362 , 11'd 1078 : cos_data <= {-16'd00143};
        11'd 363 , 11'd 1077 : cos_data <= {-16'd00214};
        11'd 364 , 11'd 1076 : cos_data <= {-16'd00286};
        11'd 365 , 11'd 1075 : cos_data <= {-16'd00357};
        11'd 366 , 11'd 1074 : cos_data <= {-16'd00429};
        11'd 367 , 11'd 1073 : cos_data <= {-16'd00500};
        11'd 368 , 11'd 1072 : cos_data <= {-16'd00572};
        11'd 369 , 11'd 1071 : cos_data <= {-16'd00643};
        11'd 370 , 11'd 1070 : cos_data <= {-16'd00715};
        11'd 371 , 11'd 1069 : cos_data <= {-16'd00786};
        11'd 372 , 11'd 1068 : cos_data <= {-16'd00857};
        11'd 373 , 11'd 1067 : cos_data <= {-16'd00929};
        11'd 374 , 11'd 1066 : cos_data <= {-16'd01000};
        11'd 375 , 11'd 1065 : cos_data <= {-16'd01072};
        11'd 376 , 11'd 1064 : cos_data <= {-16'd01143};
        11'd 377 , 11'd 1063 : cos_data <= {-16'd01214};
        11'd 378 , 11'd 1062 : cos_data <= {-16'd01285};
        11'd 379 , 11'd 1061 : cos_data <= {-16'd01357};
        11'd 380 , 11'd 1060 : cos_data <= {-16'd01428};
        11'd 381 , 11'd 1059 : cos_data <= {-16'd01499};
        11'd 382 , 11'd 1058 : cos_data <= {-16'd01570};
        11'd 383 , 11'd 1057 : cos_data <= {-16'd01641};
        11'd 384 , 11'd 1056 : cos_data <= {-16'd01713};
        11'd 385 , 11'd 1055 : cos_data <= {-16'd01784};
        11'd 386 , 11'd 1054 : cos_data <= {-16'd01855};
        11'd 387 , 11'd 1053 : cos_data <= {-16'd01926};
        11'd 388 , 11'd 1052 : cos_data <= {-16'd01997};
        11'd 389 , 11'd 1051 : cos_data <= {-16'd02068};
        11'd 390 , 11'd 1050 : cos_data <= {-16'd02139};
        11'd 391 , 11'd 1049 : cos_data <= {-16'd02209};
        11'd 392 , 11'd 1048 : cos_data <= {-16'd02280};
        11'd 393 , 11'd 1047 : cos_data <= {-16'd02351};
        11'd 394 , 11'd 1046 : cos_data <= {-16'd02422};
        11'd 395 , 11'd 1045 : cos_data <= {-16'd02492};
        11'd 396 , 11'd 1044 : cos_data <= {-16'd02563};
        11'd 397 , 11'd 1043 : cos_data <= {-16'd02634};
        11'd 398 , 11'd 1042 : cos_data <= {-16'd02704};
        11'd 399 , 11'd 1041 : cos_data <= {-16'd02775};
        11'd 400 , 11'd 1040 : cos_data <= {-16'd02845};
        11'd 401 , 11'd 1039 : cos_data <= {-16'd02915};
        11'd 402 , 11'd 1038 : cos_data <= {-16'd02986};
        11'd 403 , 11'd 1037 : cos_data <= {-16'd03056};
        11'd 404 , 11'd 1036 : cos_data <= {-16'd03126};
        11'd 405 , 11'd 1035 : cos_data <= {-16'd03196};
        11'd 406 , 11'd 1034 : cos_data <= {-16'd03266};
        11'd 407 , 11'd 1033 : cos_data <= {-16'd03336};
        11'd 408 , 11'd 1032 : cos_data <= {-16'd03406};
        11'd 409 , 11'd 1031 : cos_data <= {-16'd03476};
        11'd 410 , 11'd 1030 : cos_data <= {-16'd03546};
        11'd 411 , 11'd 1029 : cos_data <= {-16'd03616};
        11'd 412 , 11'd 1028 : cos_data <= {-16'd03686};
        11'd 413 , 11'd 1027 : cos_data <= {-16'd03755};
        11'd 414 , 11'd 1026 : cos_data <= {-16'd03825};
        11'd 415 , 11'd 1025 : cos_data <= {-16'd03894};
        11'd 416 , 11'd 1024 : cos_data <= {-16'd03964};
        11'd 417 , 11'd 1023 : cos_data <= {-16'd04033};
        11'd 418 , 11'd 1022 : cos_data <= {-16'd04102};
        11'd 419 , 11'd 1021 : cos_data <= {-16'd04171};
        11'd 420 , 11'd 1020 : cos_data <= {-16'd04240};
        11'd 421 , 11'd 1019 : cos_data <= {-16'd04310};
        11'd 422 , 11'd 1018 : cos_data <= {-16'd04378};
        11'd 423 , 11'd 1017 : cos_data <= {-16'd04447};
        11'd 424 , 11'd 1016 : cos_data <= {-16'd04516};
        11'd 425 , 11'd 1015 : cos_data <= {-16'd04585};
        11'd 426 , 11'd 1014 : cos_data <= {-16'd04653};
        11'd 427 , 11'd 1013 : cos_data <= {-16'd04722};
        11'd 428 , 11'd 1012 : cos_data <= {-16'd04790};
        11'd 429 , 11'd 1011 : cos_data <= {-16'd04859};
        11'd 430 , 11'd 1010 : cos_data <= {-16'd04927};
        11'd 431 , 11'd 1009 : cos_data <= {-16'd04995};
        11'd 432 , 11'd 1008 : cos_data <= {-16'd05063};
        11'd 433 , 11'd 1007 : cos_data <= {-16'd05131};
        11'd 434 , 11'd 1006 : cos_data <= {-16'd05199};
        11'd 435 , 11'd 1005 : cos_data <= {-16'd05266};
        11'd 436 , 11'd 1004 : cos_data <= {-16'd05334};
        11'd 437 , 11'd 1003 : cos_data <= {-16'd05402};
        11'd 438 , 11'd 1002 : cos_data <= {-16'd05469};
        11'd 439 , 11'd 1001 : cos_data <= {-16'd05536};
        11'd 440 , 11'd 1000 : cos_data <= {-16'd05604};
        11'd 441 , 11'd 999  : cos_data <= {-16'd05671};
        11'd 442 , 11'd 998  : cos_data <= {-16'd05738};
        11'd 443 , 11'd 997  : cos_data <= {-16'd05805};
        11'd 444 , 11'd 996  : cos_data <= {-16'd05872};
        11'd 445 , 11'd 995  : cos_data <= {-16'd05938};
        11'd 446 , 11'd 994  : cos_data <= {-16'd06005};
        11'd 447 , 11'd 993  : cos_data <= {-16'd06071};
        11'd 448 , 11'd 992  : cos_data <= {-16'd06138};
        11'd 449 , 11'd 991  : cos_data <= {-16'd06204};
        11'd 450 , 11'd 990  : cos_data <= {-16'd06270};
        11'd 451 , 11'd 989  : cos_data <= {-16'd06336};
        11'd 452 , 11'd 988  : cos_data <= {-16'd06402};
        11'd 453 , 11'd 987  : cos_data <= {-16'd06467};
        11'd 454 , 11'd 986  : cos_data <= {-16'd06533};
        11'd 455 , 11'd 985  : cos_data <= {-16'd06599};
        11'd 456 , 11'd 984  : cos_data <= {-16'd06664};
        11'd 457 , 11'd 983  : cos_data <= {-16'd06729};
        11'd 458 , 11'd 982  : cos_data <= {-16'd06794};
        11'd 459 , 11'd 981  : cos_data <= {-16'd06859};
        11'd 460 , 11'd 980  : cos_data <= {-16'd06924};
        11'd 461 , 11'd 979  : cos_data <= {-16'd06989};
        11'd 462 , 11'd 978  : cos_data <= {-16'd07053};
        11'd 463 , 11'd 977  : cos_data <= {-16'd07118};
        11'd 464 , 11'd 976  : cos_data <= {-16'd07182};
        11'd 465 , 11'd 975  : cos_data <= {-16'd07246};
        11'd 466 , 11'd 974  : cos_data <= {-16'd07311};
        11'd 467 , 11'd 973  : cos_data <= {-16'd07374};
        11'd 468 , 11'd 972  : cos_data <= {-16'd07438};
        11'd 469 , 11'd 971  : cos_data <= {-16'd07502};
        11'd 470 , 11'd 970  : cos_data <= {-16'd07565};
        11'd 471 , 11'd 969  : cos_data <= {-16'd07629};
        11'd 472 , 11'd 968  : cos_data <= {-16'd07692};
        11'd 473 , 11'd 967  : cos_data <= {-16'd07755};
        11'd 474 , 11'd 966  : cos_data <= {-16'd07818};
        11'd 475 , 11'd 965  : cos_data <= {-16'd07881};
        11'd 476 , 11'd 964  : cos_data <= {-16'd07943};
        11'd 477 , 11'd 963  : cos_data <= {-16'd08006};
        11'd 478 , 11'd 962  : cos_data <= {-16'd08068};
        11'd 479 , 11'd 961  : cos_data <= {-16'd08130};
        11'd 480 , 11'd 960  : cos_data <= {-16'd08192};
        11'd 481 , 11'd 959  : cos_data <= {-16'd08254};
        11'd 482 , 11'd 958  : cos_data <= {-16'd08316};
        11'd 483 , 11'd 957  : cos_data <= {-16'd08377};
        11'd 484 , 11'd 956  : cos_data <= {-16'd08438};
        11'd 485 , 11'd 955  : cos_data <= {-16'd08500};
        11'd 486 , 11'd 954  : cos_data <= {-16'd08561};
        11'd 487 , 11'd 953  : cos_data <= {-16'd08621};
        11'd 488 , 11'd 952  : cos_data <= {-16'd08682};
        11'd 489 , 11'd 951  : cos_data <= {-16'd08743};
        11'd 490 , 11'd 950  : cos_data <= {-16'd08803};
        11'd 491 , 11'd 949  : cos_data <= {-16'd08863};
        11'd 492 , 11'd 948  : cos_data <= {-16'd08923};
        11'd 493 , 11'd 947  : cos_data <= {-16'd08983};
        11'd 494 , 11'd 946  : cos_data <= {-16'd09043};
        11'd 495 , 11'd 945  : cos_data <= {-16'd09102};
        11'd 496 , 11'd 944  : cos_data <= {-16'd09162};
        11'd 497 , 11'd 943  : cos_data <= {-16'd09221};
        11'd 498 , 11'd 942  : cos_data <= {-16'd09280};
        11'd 499 , 11'd 941  : cos_data <= {-16'd09339};
        11'd 500 , 11'd 940  : cos_data <= {-16'd09397};
        11'd 501 , 11'd 939  : cos_data <= {-16'd09456};
        11'd 502 , 11'd 938  : cos_data <= {-16'd09514};
        11'd 503 , 11'd 937  : cos_data <= {-16'd09572};
        11'd 504 , 11'd 936  : cos_data <= {-16'd09630};
        11'd 505 , 11'd 935  : cos_data <= {-16'd09688};
        11'd 506 , 11'd 934  : cos_data <= {-16'd09746};
        11'd 507 , 11'd 933  : cos_data <= {-16'd09803};
        11'd 508 , 11'd 932  : cos_data <= {-16'd09860};
        11'd 509 , 11'd 931  : cos_data <= {-16'd09917};
        11'd 510 , 11'd 930  : cos_data <= {-16'd09974};
        11'd 511 , 11'd 929  : cos_data <= {-16'd10031};
        11'd 512 , 11'd 928  : cos_data <= {-16'd10087};
        11'd 513 , 11'd 927  : cos_data <= {-16'd10143};
        11'd 514 , 11'd 926  : cos_data <= {-16'd10199};
        11'd 515 , 11'd 925  : cos_data <= {-16'd10255};
        11'd 516 , 11'd 924  : cos_data <= {-16'd10311};
        11'd 517 , 11'd 923  : cos_data <= {-16'd10366};
        11'd 518 , 11'd 922  : cos_data <= {-16'd10422};
        11'd 519 , 11'd 921  : cos_data <= {-16'd10477};
        11'd 520 , 11'd 920  : cos_data <= {-16'd10531};
        11'd 521 , 11'd 919  : cos_data <= {-16'd10586};
        11'd 522 , 11'd 918  : cos_data <= {-16'd10641};
        11'd 523 , 11'd 917  : cos_data <= {-16'd10695};
        11'd 524 , 11'd 916  : cos_data <= {-16'd10749};
        11'd 525 , 11'd 915  : cos_data <= {-16'd10803};
        11'd 526 , 11'd 914  : cos_data <= {-16'd10856};
        11'd 527 , 11'd 913  : cos_data <= {-16'd10910};
        11'd 528 , 11'd 912  : cos_data <= {-16'd10963};
        11'd 529 , 11'd 911  : cos_data <= {-16'd11016};
        11'd 530 , 11'd 910  : cos_data <= {-16'd11069};
        11'd 531 , 11'd 909  : cos_data <= {-16'd11121};
        11'd 532 , 11'd 908  : cos_data <= {-16'd11174};
        11'd 533 , 11'd 907  : cos_data <= {-16'd11226};
        11'd 534 , 11'd 906  : cos_data <= {-16'd11278};
        11'd 535 , 11'd 905  : cos_data <= {-16'd11330};
        11'd 536 , 11'd 904  : cos_data <= {-16'd11381};
        11'd 537 , 11'd 903  : cos_data <= {-16'd11433};
        11'd 538 , 11'd 902  : cos_data <= {-16'd11484};
        11'd 539 , 11'd 901  : cos_data <= {-16'd11535};
        11'd 540 , 11'd 900  : cos_data <= {-16'd11585};
        11'd 541 , 11'd 899  : cos_data <= {-16'd11636};
        11'd 542 , 11'd 898  : cos_data <= {-16'd11686};
        11'd 543 , 11'd 897  : cos_data <= {-16'd11736};
        11'd 544 , 11'd 896  : cos_data <= {-16'd11786};
        11'd 545 , 11'd 895  : cos_data <= {-16'd11835};
        11'd 546 , 11'd 894  : cos_data <= {-16'd11885};
        11'd 547 , 11'd 893  : cos_data <= {-16'd11934};
        11'd 548 , 11'd 892  : cos_data <= {-16'd11982};
        11'd 549 , 11'd 891  : cos_data <= {-16'd12031};
        11'd 550 , 11'd 890  : cos_data <= {-16'd12080};
        11'd 551 , 11'd 889  : cos_data <= {-16'd12128};
        11'd 552 , 11'd 888  : cos_data <= {-16'd12176};
        11'd 553 , 11'd 887  : cos_data <= {-16'd12223};
        11'd 554 , 11'd 886  : cos_data <= {-16'd12271};
        11'd 555 , 11'd 885  : cos_data <= {-16'd12318};
        11'd 556 , 11'd 884  : cos_data <= {-16'd12365};
        11'd 557 , 11'd 883  : cos_data <= {-16'd12412};
        11'd 558 , 11'd 882  : cos_data <= {-16'd12458};
        11'd 559 , 11'd 881  : cos_data <= {-16'd12505};
        11'd 560 , 11'd 880  : cos_data <= {-16'd12551};
        11'd 561 , 11'd 879  : cos_data <= {-16'd12597};
        11'd 562 , 11'd 878  : cos_data <= {-16'd12642};
        11'd 563 , 11'd 877  : cos_data <= {-16'd12688};
        11'd 564 , 11'd 876  : cos_data <= {-16'd12733};
        11'd 565 , 11'd 875  : cos_data <= {-16'd12778};
        11'd 566 , 11'd 874  : cos_data <= {-16'd12822};
        11'd 567 , 11'd 873  : cos_data <= {-16'd12867};
        11'd 568 , 11'd 872  : cos_data <= {-16'd12911};
        11'd 569 , 11'd 871  : cos_data <= {-16'd12955};
        11'd 570 , 11'd 870  : cos_data <= {-16'd12998};
        11'd 571 , 11'd 869  : cos_data <= {-16'd13042};
        11'd 572 , 11'd 868  : cos_data <= {-16'd13085};
        11'd 573 , 11'd 867  : cos_data <= {-16'd13128};
        11'd 574 , 11'd 866  : cos_data <= {-16'd13170};
        11'd 575 , 11'd 865  : cos_data <= {-16'd13213};
        11'd 576 , 11'd 864  : cos_data <= {-16'd13255};
        11'd 577 , 11'd 863  : cos_data <= {-16'd13297};
        11'd 578 , 11'd 862  : cos_data <= {-16'd13338};
        11'd 579 , 11'd 861  : cos_data <= {-16'd13380};
        11'd 580 , 11'd 860  : cos_data <= {-16'd13421};
        11'd 581 , 11'd 859  : cos_data <= {-16'd13462};
        11'd 582 , 11'd 858  : cos_data <= {-16'd13502};
        11'd 583 , 11'd 857  : cos_data <= {-16'd13543};
        11'd 584 , 11'd 856  : cos_data <= {-16'd13583};
        11'd 585 , 11'd 855  : cos_data <= {-16'd13623};
        11'd 586 , 11'd 854  : cos_data <= {-16'd13662};
        11'd 587 , 11'd 853  : cos_data <= {-16'd13702};
        11'd 588 , 11'd 852  : cos_data <= {-16'd13741};
        11'd 589 , 11'd 851  : cos_data <= {-16'd13780};
        11'd 590 , 11'd 850  : cos_data <= {-16'd13818};
        11'd 591 , 11'd 849  : cos_data <= {-16'd13856};
        11'd 592 , 11'd 848  : cos_data <= {-16'd13894};
        11'd 593 , 11'd 847  : cos_data <= {-16'd13932};
        11'd 594 , 11'd 846  : cos_data <= {-16'd13970};
        11'd 595 , 11'd 845  : cos_data <= {-16'd14007};
        11'd 596 , 11'd 844  : cos_data <= {-16'd14044};
        11'd 597 , 11'd 843  : cos_data <= {-16'd14081};
        11'd 598 , 11'd 842  : cos_data <= {-16'd14117};
        11'd 599 , 11'd 841  : cos_data <= {-16'd14153};
        11'd 600 , 11'd 840  : cos_data <= {-16'd14189};
        11'd 601 , 11'd 839  : cos_data <= {-16'd14225};
        11'd 602 , 11'd 838  : cos_data <= {-16'd14260};
        11'd 603 , 11'd 837  : cos_data <= {-16'd14295};
        11'd 604 , 11'd 836  : cos_data <= {-16'd14330};
        11'd 605 , 11'd 835  : cos_data <= {-16'd14364};
        11'd 606 , 11'd 834  : cos_data <= {-16'd14399};
        11'd 607 , 11'd 833  : cos_data <= {-16'd14433};
        11'd 608 , 11'd 832  : cos_data <= {-16'd14466};
        11'd 609 , 11'd 831  : cos_data <= {-16'd14500};
        11'd 610 , 11'd 830  : cos_data <= {-16'd14533};
        11'd 611 , 11'd 829  : cos_data <= {-16'd14566};
        11'd 612 , 11'd 828  : cos_data <= {-16'd14598};
        11'd 613 , 11'd 827  : cos_data <= {-16'd14631};
        11'd 614 , 11'd 826  : cos_data <= {-16'd14663};
        11'd 615 , 11'd 825  : cos_data <= {-16'd14694};
        11'd 616 , 11'd 824  : cos_data <= {-16'd14726};
        11'd 617 , 11'd 823  : cos_data <= {-16'd14757};
        11'd 618 , 11'd 822  : cos_data <= {-16'd14788};
        11'd 619 , 11'd 821  : cos_data <= {-16'd14819};
        11'd 620 , 11'd 820  : cos_data <= {-16'd14849};
        11'd 621 , 11'd 819  : cos_data <= {-16'd14879};
        11'd 622 , 11'd 818  : cos_data <= {-16'd14909};
        11'd 623 , 11'd 817  : cos_data <= {-16'd14938};
        11'd 624 , 11'd 816  : cos_data <= {-16'd14968};
        11'd 625 , 11'd 815  : cos_data <= {-16'd14996};
        11'd 626 , 11'd 814  : cos_data <= {-16'd15025};
        11'd 627 , 11'd 813  : cos_data <= {-16'd15053};
        11'd 628 , 11'd 812  : cos_data <= {-16'd15082};
        11'd 629 , 11'd 811  : cos_data <= {-16'd15109};
        11'd 630 , 11'd 810  : cos_data <= {-16'd15137};
        11'd 631 , 11'd 809  : cos_data <= {-16'd15164};
        11'd 632 , 11'd 808  : cos_data <= {-16'd15191};
        11'd 633 , 11'd 807  : cos_data <= {-16'd15218};
        11'd 634 , 11'd 806  : cos_data <= {-16'd15244};
        11'd 635 , 11'd 805  : cos_data <= {-16'd15270};
        11'd 636 , 11'd 804  : cos_data <= {-16'd15296};
        11'd 637 , 11'd 803  : cos_data <= {-16'd15321};
        11'd 638 , 11'd 802  : cos_data <= {-16'd15346};
        11'd 639 , 11'd 801  : cos_data <= {-16'd15371};
        11'd 640 , 11'd 800  : cos_data <= {-16'd15396};
        11'd 641 , 11'd 799  : cos_data <= {-16'd15420};
        11'd 642 , 11'd 798  : cos_data <= {-16'd15444};
        11'd 643 , 11'd 797  : cos_data <= {-16'd15468};
        11'd 644 , 11'd 796  : cos_data <= {-16'd15491};
        11'd 645 , 11'd 795  : cos_data <= {-16'd15515};
        11'd 646 , 11'd 794  : cos_data <= {-16'd15537};
        11'd 647 , 11'd 793  : cos_data <= {-16'd15560};
        11'd 648 , 11'd 792  : cos_data <= {-16'd15582};
        11'd 649 , 11'd 791  : cos_data <= {-16'd15604};
        11'd 650 , 11'd 790  : cos_data <= {-16'd15626};
        11'd 651 , 11'd 789  : cos_data <= {-16'd15647};
        11'd 652 , 11'd 788  : cos_data <= {-16'd15668};
        11'd 653 , 11'd 787  : cos_data <= {-16'd15689};
        11'd 654 , 11'd 786  : cos_data <= {-16'd15709};
        11'd 655 , 11'd 785  : cos_data <= {-16'd15729};
        11'd 656 , 11'd 784  : cos_data <= {-16'd15749};
        11'd 657 , 11'd 783  : cos_data <= {-16'd15769};
        11'd 658 , 11'd 782  : cos_data <= {-16'd15788};
        11'd 659 , 11'd 781  : cos_data <= {-16'd15807};
        11'd 660 , 11'd 780  : cos_data <= {-16'd15826};
        11'd 661 , 11'd 779  : cos_data <= {-16'd15844};
        11'd 662 , 11'd 778  : cos_data <= {-16'd15862};
        11'd 663 , 11'd 777  : cos_data <= {-16'd15880};
        11'd 664 , 11'd 776  : cos_data <= {-16'd15897};
        11'd 665 , 11'd 775  : cos_data <= {-16'd15914};
        11'd 666 , 11'd 774  : cos_data <= {-16'd15931};
        11'd 667 , 11'd 773  : cos_data <= {-16'd15948};
        11'd 668 , 11'd 772  : cos_data <= {-16'd15964};
        11'd 669 , 11'd 771  : cos_data <= {-16'd15980};
        11'd 670 , 11'd 770  : cos_data <= {-16'd15996};
        11'd 671 , 11'd 769  : cos_data <= {-16'd16011};
        11'd 672 , 11'd 768  : cos_data <= {-16'd16026};
        11'd 673 , 11'd 767  : cos_data <= {-16'd16041};
        11'd 674 , 11'd 766  : cos_data <= {-16'd16055};
        11'd 675 , 11'd 765  : cos_data <= {-16'd16069};
        11'd 676 , 11'd 764  : cos_data <= {-16'd16083};
        11'd 677 , 11'd 763  : cos_data <= {-16'd16096};
        11'd 678 , 11'd 762  : cos_data <= {-16'd16110};
        11'd 679 , 11'd 761  : cos_data <= {-16'd16123};
        11'd 680 , 11'd 760  : cos_data <= {-16'd16135};
        11'd 681 , 11'd 759  : cos_data <= {-16'd16147};
        11'd 682 , 11'd 758  : cos_data <= {-16'd16159};
        11'd 683 , 11'd 757  : cos_data <= {-16'd16171};
        11'd 684 , 11'd 756  : cos_data <= {-16'd16182};
        11'd 685 , 11'd 755  : cos_data <= {-16'd16193};
        11'd 686 , 11'd 754  : cos_data <= {-16'd16204};
        11'd 687 , 11'd 753  : cos_data <= {-16'd16214};
        11'd 688 , 11'd 752  : cos_data <= {-16'd16225};
        11'd 689 , 11'd 751  : cos_data <= {-16'd16234};
        11'd 690 , 11'd 750  : cos_data <= {-16'd16244};
        11'd 691 , 11'd 749  : cos_data <= {-16'd16253};
        11'd 692 , 11'd 748  : cos_data <= {-16'd16262};
        11'd 693 , 11'd 747  : cos_data <= {-16'd16270};
        11'd 694 , 11'd 746  : cos_data <= {-16'd16279};
        11'd 695 , 11'd 745  : cos_data <= {-16'd16287};
        11'd 696 , 11'd 744  : cos_data <= {-16'd16294};
        11'd 697 , 11'd 743  : cos_data <= {-16'd16302};
        11'd 698 , 11'd 742  : cos_data <= {-16'd16309};
        11'd 699 , 11'd 741  : cos_data <= {-16'd16315};
        11'd 700 , 11'd 740  : cos_data <= {-16'd16322};
        11'd 701 , 11'd 739  : cos_data <= {-16'd16328};
        11'd 702 , 11'd 738  : cos_data <= {-16'd16333};
        11'd 703 , 11'd 737  : cos_data <= {-16'd16339};
        11'd 704 , 11'd 736  : cos_data <= {-16'd16344};
        11'd 705 , 11'd 735  : cos_data <= {-16'd16349};
        11'd 706 , 11'd 734  : cos_data <= {-16'd16353};
        11'd 707 , 11'd 733  : cos_data <= {-16'd16358};
        11'd 708 , 11'd 732  : cos_data <= {-16'd16362};
        11'd 709 , 11'd 731  : cos_data <= {-16'd16365};
        11'd 710 , 11'd 730  : cos_data <= {-16'd16368};
        11'd 711 , 11'd 729  : cos_data <= {-16'd16371};
        11'd 712 , 11'd 728  : cos_data <= {-16'd16374};
        11'd 713 , 11'd 727  : cos_data <= {-16'd16376};
        11'd 714 , 11'd 726  : cos_data <= {-16'd16378};
        11'd 715 , 11'd 725  : cos_data <= {-16'd16380};
        11'd 716 , 11'd 724  : cos_data <= {-16'd16382};
        11'd 717 , 11'd 723  : cos_data <= {-16'd16383};
        11'd 718 , 11'd 722  : cos_data <= {-16'd16383};
        11'd 719 , 11'd 721  : cos_data <= {-16'd16384};
        11'd 720             : cos_data <= {-16'd16384};
        
        default: cos_data <= {16'd16384};
    endcase
end

endmodule

