module lut_4sin16384(
    input[9:0]             lut_index,
    output reg[31:0]       lut_data
);

always@(*) begin
    case(lut_index)
        10'd    1: lut_data <= {10'd00071};
        10'd    2: lut_data <= {10'd00143};
        10'd    3: lut_data <= {10'd00214};
        10'd    4: lut_data <= {10'd00286};
        10'd    5: lut_data <= {10'd00357};
        10'd    6: lut_data <= {10'd00429};
        10'd    7: lut_data <= {10'd00500};
        10'd    8: lut_data <= {10'd00572};
        10'd    9: lut_data <= {10'd00643};
        10'd   10: lut_data <= {10'd00715};
        10'd   11: lut_data <= {10'd00786};
        10'd   12: lut_data <= {10'd00857};
        10'd   13: lut_data <= {10'd00929};
        10'd   14: lut_data <= {10'd01000};
        10'd   15: lut_data <= {10'd01072};
        10'd   16: lut_data <= {10'd01143};
        10'd   17: lut_data <= {10'd01214};
        10'd   18: lut_data <= {10'd01285};
        10'd   19: lut_data <= {10'd01357};
        10'd   20: lut_data <= {10'd01428};
        10'd   21: lut_data <= {10'd01499};
        10'd   22: lut_data <= {10'd01570};
        10'd   23: lut_data <= {10'd01641};
        10'd   24: lut_data <= {10'd01713};
        10'd   25: lut_data <= {10'd01784};
        10'd   26: lut_data <= {10'd01855};
        10'd   27: lut_data <= {10'd01926};
        10'd   28: lut_data <= {10'd01997};
        10'd   29: lut_data <= {10'd02068};
        10'd   30: lut_data <= {10'd02139};
        10'd   31: lut_data <= {10'd02209};
        10'd   32: lut_data <= {10'd02280};
        10'd   33: lut_data <= {10'd02351};
        10'd   34: lut_data <= {10'd02422};
        10'd   35: lut_data <= {10'd02492};
        10'd   36: lut_data <= {10'd02563};
        10'd   37: lut_data <= {10'd02634};
        10'd   38: lut_data <= {10'd02704};
        10'd   39: lut_data <= {10'd02775};
        10'd   40: lut_data <= {10'd02845};
        10'd   41: lut_data <= {10'd02915};
        10'd   42: lut_data <= {10'd02986};
        10'd   43: lut_data <= {10'd03056};
        10'd   44: lut_data <= {10'd03126};
        10'd   45: lut_data <= {10'd03196};
        10'd   46: lut_data <= {10'd03266};
        10'd   47: lut_data <= {10'd03336};
        10'd   48: lut_data <= {10'd03406};
        10'd   49: lut_data <= {10'd03476};
        10'd   50: lut_data <= {10'd03546};
        10'd   51: lut_data <= {10'd03616};
        10'd   52: lut_data <= {10'd03686};
        10'd   53: lut_data <= {10'd03755};
        10'd   54: lut_data <= {10'd03825};
        10'd   55: lut_data <= {10'd03894};
        10'd   56: lut_data <= {10'd03964};
        10'd   57: lut_data <= {10'd04033};
        10'd   58: lut_data <= {10'd04102};
        10'd   59: lut_data <= {10'd04171};
        10'd   60: lut_data <= {10'd04240};
        10'd   61: lut_data <= {10'd04310};
        10'd   62: lut_data <= {10'd04378};
        10'd   63: lut_data <= {10'd04447};
        10'd   64: lut_data <= {10'd04516};
        10'd   65: lut_data <= {10'd04585};
        10'd   66: lut_data <= {10'd04653};
        10'd   67: lut_data <= {10'd04722};
        10'd   68: lut_data <= {10'd04790};
        10'd   69: lut_data <= {10'd04859};
        10'd   70: lut_data <= {10'd04927};
        10'd   71: lut_data <= {10'd04995};
        10'd   72: lut_data <= {10'd05063};
        10'd   73: lut_data <= {10'd05131};
        10'd   74: lut_data <= {10'd05199};
        10'd   75: lut_data <= {10'd05266};
        10'd   76: lut_data <= {10'd05334};
        10'd   77: lut_data <= {10'd05402};
        10'd   78: lut_data <= {10'd05469};
        10'd   79: lut_data <= {10'd05536};
        10'd   80: lut_data <= {10'd05604};
        10'd   81: lut_data <= {10'd05671};
        10'd   82: lut_data <= {10'd05738};
        10'd   83: lut_data <= {10'd05805};
        10'd   84: lut_data <= {10'd05872};
        10'd   85: lut_data <= {10'd05938};
        10'd   86: lut_data <= {10'd06005};
        10'd   87: lut_data <= {10'd06071};
        10'd   88: lut_data <= {10'd06138};
        10'd   89: lut_data <= {10'd06204};
        10'd   90: lut_data <= {10'd06270};
        10'd   91: lut_data <= {10'd06336};
        10'd   92: lut_data <= {10'd06402};
        10'd   93: lut_data <= {10'd06467};
        10'd   94: lut_data <= {10'd06533};
        10'd   95: lut_data <= {10'd06599};
        10'd   96: lut_data <= {10'd06664};
        10'd   97: lut_data <= {10'd06729};
        10'd   98: lut_data <= {10'd06794};
        10'd   99: lut_data <= {10'd06859};
        10'd  100: lut_data <= {10'd06924};
        10'd  101: lut_data <= {10'd06989};
        10'd  102: lut_data <= {10'd07053};
        10'd  103: lut_data <= {10'd07118};
        10'd  104: lut_data <= {10'd07182};
        10'd  105: lut_data <= {10'd07246};
        10'd  106: lut_data <= {10'd07311};
        10'd  107: lut_data <= {10'd07374};
        10'd  108: lut_data <= {10'd07438};
        10'd  109: lut_data <= {10'd07502};
        10'd  110: lut_data <= {10'd07565};
        10'd  111: lut_data <= {10'd07629};
        10'd  112: lut_data <= {10'd07692};
        10'd  113: lut_data <= {10'd07755};
        10'd  114: lut_data <= {10'd07818};
        10'd  115: lut_data <= {10'd07881};
        10'd  116: lut_data <= {10'd07943};
        10'd  117: lut_data <= {10'd08006};
        10'd  118: lut_data <= {10'd08068};
        10'd  119: lut_data <= {10'd08130};
        10'd  120: lut_data <= {10'd08192};
        10'd  121: lut_data <= {10'd08254};
        10'd  122: lut_data <= {10'd08316};
        10'd  123: lut_data <= {10'd08377};
        10'd  124: lut_data <= {10'd08438};
        10'd  125: lut_data <= {10'd08500};
        10'd  126: lut_data <= {10'd08561};
        10'd  127: lut_data <= {10'd08621};
        10'd  128: lut_data <= {10'd08682};
        10'd  129: lut_data <= {10'd08743};
        10'd  130: lut_data <= {10'd08803};
        10'd  131: lut_data <= {10'd08863};
        10'd  132: lut_data <= {10'd08923};
        10'd  133: lut_data <= {10'd08983};
        10'd  134: lut_data <= {10'd09043};
        10'd  135: lut_data <= {10'd09102};
        10'd  136: lut_data <= {10'd09162};
        10'd  137: lut_data <= {10'd09221};
        10'd  138: lut_data <= {10'd09280};
        10'd  139: lut_data <= {10'd09339};
        10'd  140: lut_data <= {10'd09397};
        10'd  141: lut_data <= {10'd09456};
        10'd  142: lut_data <= {10'd09514};
        10'd  143: lut_data <= {10'd09572};
        10'd  144: lut_data <= {10'd09630};
        10'd  145: lut_data <= {10'd09688};
        10'd  146: lut_data <= {10'd09746};
        10'd  147: lut_data <= {10'd09803};
        10'd  148: lut_data <= {10'd09860};
        10'd  149: lut_data <= {10'd09917};
        10'd  150: lut_data <= {10'd09974};
        10'd  151: lut_data <= {10'd10031};
        10'd  152: lut_data <= {10'd10087};
        10'd  153: lut_data <= {10'd10143};
        10'd  154: lut_data <= {10'd10199};
        10'd  155: lut_data <= {10'd10255};
        10'd  156: lut_data <= {10'd10311};
        10'd  157: lut_data <= {10'd10366};
        10'd  158: lut_data <= {10'd10422};
        10'd  159: lut_data <= {10'd10477};
        10'd  160: lut_data <= {10'd10531};
        10'd  161: lut_data <= {10'd10586};
        10'd  162: lut_data <= {10'd10641};
        10'd  163: lut_data <= {10'd10695};
        10'd  164: lut_data <= {10'd10749};
        10'd  165: lut_data <= {10'd10803};
        10'd  166: lut_data <= {10'd10856};
        10'd  167: lut_data <= {10'd10910};
        10'd  168: lut_data <= {10'd10963};
        10'd  169: lut_data <= {10'd11016};
        10'd  170: lut_data <= {10'd11069};
        10'd  171: lut_data <= {10'd11121};
        10'd  172: lut_data <= {10'd11174};
        10'd  173: lut_data <= {10'd11226};
        10'd  174: lut_data <= {10'd11278};
        10'd  175: lut_data <= {10'd11330};
        10'd  176: lut_data <= {10'd11381};
        10'd  177: lut_data <= {10'd11433};
        10'd  178: lut_data <= {10'd11484};
        10'd  179: lut_data <= {10'd11535};
        10'd  180: lut_data <= {10'd11585};
        10'd  181: lut_data <= {10'd11636};
        10'd  182: lut_data <= {10'd11686};
        10'd  183: lut_data <= {10'd11736};
        10'd  184: lut_data <= {10'd11786};
        10'd  185: lut_data <= {10'd11835};
        10'd  186: lut_data <= {10'd11885};
        10'd  187: lut_data <= {10'd11934};
        10'd  188: lut_data <= {10'd11982};
        10'd  189: lut_data <= {10'd12031};
        10'd  190: lut_data <= {10'd12080};
        10'd  191: lut_data <= {10'd12128};
        10'd  192: lut_data <= {10'd12176};
        10'd  193: lut_data <= {10'd12223};
        10'd  194: lut_data <= {10'd12271};
        10'd  195: lut_data <= {10'd12318};
        10'd  196: lut_data <= {10'd12365};
        10'd  197: lut_data <= {10'd12412};
        10'd  198: lut_data <= {10'd12458};
        10'd  199: lut_data <= {10'd12505};
        10'd  200: lut_data <= {10'd12551};
        10'd  201: lut_data <= {10'd12597};
        10'd  202: lut_data <= {10'd12642};
        10'd  203: lut_data <= {10'd12688};
        10'd  204: lut_data <= {10'd12733};
        10'd  205: lut_data <= {10'd12778};
        10'd  206: lut_data <= {10'd12822};
        10'd  207: lut_data <= {10'd12867};
        10'd  208: lut_data <= {10'd12911};
        10'd  209: lut_data <= {10'd12955};
        10'd  210: lut_data <= {10'd12998};
        10'd  211: lut_data <= {10'd13042};
        10'd  212: lut_data <= {10'd13085};
        10'd  213: lut_data <= {10'd13128};
        10'd  214: lut_data <= {10'd13170};
        10'd  215: lut_data <= {10'd13213};
        10'd  216: lut_data <= {10'd13255};
        10'd  217: lut_data <= {10'd13297};
        10'd  218: lut_data <= {10'd13338};
        10'd  219: lut_data <= {10'd13380};
        10'd  220: lut_data <= {10'd13421};
        10'd  221: lut_data <= {10'd13462};
        10'd  222: lut_data <= {10'd13502};
        10'd  223: lut_data <= {10'd13543};
        10'd  224: lut_data <= {10'd13583};
        10'd  225: lut_data <= {10'd13623};
        10'd  226: lut_data <= {10'd13662};
        10'd  227: lut_data <= {10'd13702};
        10'd  228: lut_data <= {10'd13741};
        10'd  229: lut_data <= {10'd13780};
        10'd  230: lut_data <= {10'd13818};
        10'd  231: lut_data <= {10'd13856};
        10'd  232: lut_data <= {10'd13894};
        10'd  233: lut_data <= {10'd13932};
        10'd  234: lut_data <= {10'd13970};
        10'd  235: lut_data <= {10'd14007};
        10'd  236: lut_data <= {10'd14044};
        10'd  237: lut_data <= {10'd14081};
        10'd  238: lut_data <= {10'd14117};
        10'd  239: lut_data <= {10'd14153};
        10'd  240: lut_data <= {10'd14189};
        10'd  241: lut_data <= {10'd14225};
        10'd  242: lut_data <= {10'd14260};
        10'd  243: lut_data <= {10'd14295};
        10'd  244: lut_data <= {10'd14330};
        10'd  245: lut_data <= {10'd14364};
        10'd  246: lut_data <= {10'd14399};
        10'd  247: lut_data <= {10'd14433};
        10'd  248: lut_data <= {10'd14466};
        10'd  249: lut_data <= {10'd14500};
        10'd  250: lut_data <= {10'd14533};
        10'd  251: lut_data <= {10'd14566};
        10'd  252: lut_data <= {10'd14598};
        10'd  253: lut_data <= {10'd14631};
        10'd  254: lut_data <= {10'd14663};
        10'd  255: lut_data <= {10'd14694};
        10'd  256: lut_data <= {10'd14726};
        10'd  257: lut_data <= {10'd14757};
        10'd  258: lut_data <= {10'd14788};
        10'd  259: lut_data <= {10'd14819};
        10'd  260: lut_data <= {10'd14849};
        10'd  261: lut_data <= {10'd14879};
        10'd  262: lut_data <= {10'd14909};
        10'd  263: lut_data <= {10'd14938};
        10'd  264: lut_data <= {10'd14968};
        10'd  265: lut_data <= {10'd14996};
        10'd  266: lut_data <= {10'd15025};
        10'd  267: lut_data <= {10'd15053};
        10'd  268: lut_data <= {10'd15082};
        10'd  269: lut_data <= {10'd15109};
        10'd  270: lut_data <= {10'd15137};
        10'd  271: lut_data <= {10'd15164};
        10'd  272: lut_data <= {10'd15191};
        10'd  273: lut_data <= {10'd15218};
        10'd  274: lut_data <= {10'd15244};
        10'd  275: lut_data <= {10'd15270};
        10'd  276: lut_data <= {10'd15296};
        10'd  277: lut_data <= {10'd15321};
        10'd  278: lut_data <= {10'd15346};
        10'd  279: lut_data <= {10'd15371};
        10'd  280: lut_data <= {10'd15396};
        10'd  281: lut_data <= {10'd15420};
        10'd  282: lut_data <= {10'd15444};
        10'd  283: lut_data <= {10'd15468};
        10'd  284: lut_data <= {10'd15491};
        10'd  285: lut_data <= {10'd15515};
        10'd  286: lut_data <= {10'd15537};
        10'd  287: lut_data <= {10'd15560};
        10'd  288: lut_data <= {10'd15582};
        10'd  289: lut_data <= {10'd15604};
        10'd  290: lut_data <= {10'd15626};
        10'd  291: lut_data <= {10'd15647};
        10'd  292: lut_data <= {10'd15668};
        10'd  293: lut_data <= {10'd15689};
        10'd  294: lut_data <= {10'd15709};
        10'd  295: lut_data <= {10'd15729};
        10'd  296: lut_data <= {10'd15749};
        10'd  297: lut_data <= {10'd15769};
        10'd  298: lut_data <= {10'd15788};
        10'd  299: lut_data <= {10'd15807};
        10'd  300: lut_data <= {10'd15826};
        10'd  301: lut_data <= {10'd15844};
        10'd  302: lut_data <= {10'd15862};
        10'd  303: lut_data <= {10'd15880};
        10'd  304: lut_data <= {10'd15897};
        10'd  305: lut_data <= {10'd15914};
        10'd  306: lut_data <= {10'd15931};
        10'd  307: lut_data <= {10'd15948};
        10'd  308: lut_data <= {10'd15964};
        10'd  309: lut_data <= {10'd15980};
        10'd  310: lut_data <= {10'd15996};
        10'd  311: lut_data <= {10'd16011};
        10'd  312: lut_data <= {10'd16026};
        10'd  313: lut_data <= {10'd16041};
        10'd  314: lut_data <= {10'd16055};
        10'd  315: lut_data <= {10'd16069};
        10'd  316: lut_data <= {10'd16083};
        10'd  317: lut_data <= {10'd16096};
        10'd  318: lut_data <= {10'd16110};
        10'd  319: lut_data <= {10'd16123};
        10'd  320: lut_data <= {10'd16135};
        10'd  321: lut_data <= {10'd16147};
        10'd  322: lut_data <= {10'd16159};
        10'd  323: lut_data <= {10'd16171};
        10'd  324: lut_data <= {10'd16182};
        10'd  325: lut_data <= {10'd16193};
        10'd  326: lut_data <= {10'd16204};
        10'd  327: lut_data <= {10'd16214};
        10'd  328: lut_data <= {10'd16225};
        10'd  329: lut_data <= {10'd16234};
        10'd  330: lut_data <= {10'd16244};
        10'd  331: lut_data <= {10'd16253};
        10'd  332: lut_data <= {10'd16262};
        10'd  333: lut_data <= {10'd16270};
        10'd  334: lut_data <= {10'd16279};
        10'd  335: lut_data <= {10'd16287};
        10'd  336: lut_data <= {10'd16294};
        10'd  337: lut_data <= {10'd16302};
        10'd  338: lut_data <= {10'd16309};
        10'd  339: lut_data <= {10'd16315};
        10'd  340: lut_data <= {10'd16322};
        10'd  341: lut_data <= {10'd16328};
        10'd  342: lut_data <= {10'd16333};
        10'd  343: lut_data <= {10'd16339};
        10'd  344: lut_data <= {10'd16344};
        10'd  345: lut_data <= {10'd16349};
        10'd  346: lut_data <= {10'd16353};
        10'd  347: lut_data <= {10'd16358};
        10'd  348: lut_data <= {10'd16362};
        10'd  349: lut_data <= {10'd16365};
        10'd  350: lut_data <= {10'd16368};
        10'd  351: lut_data <= {10'd16371};
        10'd  352: lut_data <= {10'd16374};
        10'd  353: lut_data <= {10'd16376};
        10'd  354: lut_data <= {10'd16378};
        10'd  355: lut_data <= {10'd16380};
        10'd  356: lut_data <= {10'd16382};
        10'd  357: lut_data <= {10'd16383};
        10'd  358: lut_data <= {10'd16383};
        10'd  359: lut_data <= {10'd16384};
        10'd  360: lut_data <= {10'd16384};
        10'd  361: lut_data <= {10'd16384};
        10'd  362: lut_data <= {10'd16383};
        10'd  363: lut_data <= {10'd16383};
        10'd  364: lut_data <= {10'd16382};
        10'd  365: lut_data <= {10'd16380};
        10'd  366: lut_data <= {10'd16378};
        10'd  367: lut_data <= {10'd16376};
        10'd  368: lut_data <= {10'd16374};
        10'd  369: lut_data <= {10'd16371};
        10'd  370: lut_data <= {10'd16368};
        10'd  371: lut_data <= {10'd16365};
        10'd  372: lut_data <= {10'd16362};
        10'd  373: lut_data <= {10'd16358};
        10'd  374: lut_data <= {10'd16353};
        10'd  375: lut_data <= {10'd16349};
        10'd  376: lut_data <= {10'd16344};
        10'd  377: lut_data <= {10'd16339};
        10'd  378: lut_data <= {10'd16333};
        10'd  379: lut_data <= {10'd16328};
        10'd  380: lut_data <= {10'd16322};
        10'd  381: lut_data <= {10'd16315};
        10'd  382: lut_data <= {10'd16309};
        10'd  383: lut_data <= {10'd16302};
        10'd  384: lut_data <= {10'd16294};
        10'd  385: lut_data <= {10'd16287};
        10'd  386: lut_data <= {10'd16279};
        10'd  387: lut_data <= {10'd16270};
        10'd  388: lut_data <= {10'd16262};
        10'd  389: lut_data <= {10'd16253};
        10'd  390: lut_data <= {10'd16244};
        10'd  391: lut_data <= {10'd16234};
        10'd  392: lut_data <= {10'd16225};
        10'd  393: lut_data <= {10'd16214};
        10'd  394: lut_data <= {10'd16204};
        10'd  395: lut_data <= {10'd16193};
        10'd  396: lut_data <= {10'd16182};
        10'd  397: lut_data <= {10'd16171};
        10'd  398: lut_data <= {10'd16159};
        10'd  399: lut_data <= {10'd16147};
        10'd  400: lut_data <= {10'd16135};
        10'd  401: lut_data <= {10'd16123};
        10'd  402: lut_data <= {10'd16110};
        10'd  403: lut_data <= {10'd16096};
        10'd  404: lut_data <= {10'd16083};
        10'd  405: lut_data <= {10'd16069};
        10'd  406: lut_data <= {10'd16055};
        10'd  407: lut_data <= {10'd16041};
        10'd  408: lut_data <= {10'd16026};
        10'd  409: lut_data <= {10'd16011};
        10'd  410: lut_data <= {10'd15996};
        10'd  411: lut_data <= {10'd15980};
        10'd  412: lut_data <= {10'd15964};
        10'd  413: lut_data <= {10'd15948};
        10'd  414: lut_data <= {10'd15931};
        10'd  415: lut_data <= {10'd15914};
        10'd  416: lut_data <= {10'd15897};
        10'd  417: lut_data <= {10'd15880};
        10'd  418: lut_data <= {10'd15862};
        10'd  419: lut_data <= {10'd15844};
        10'd  420: lut_data <= {10'd15826};
        10'd  421: lut_data <= {10'd15807};
        10'd  422: lut_data <= {10'd15788};
        10'd  423: lut_data <= {10'd15769};
        10'd  424: lut_data <= {10'd15749};
        10'd  425: lut_data <= {10'd15729};
        10'd  426: lut_data <= {10'd15709};
        10'd  427: lut_data <= {10'd15689};
        10'd  428: lut_data <= {10'd15668};
        10'd  429: lut_data <= {10'd15647};
        10'd  430: lut_data <= {10'd15626};
        10'd  431: lut_data <= {10'd15604};
        10'd  432: lut_data <= {10'd15582};
        10'd  433: lut_data <= {10'd15560};
        10'd  434: lut_data <= {10'd15537};
        10'd  435: lut_data <= {10'd15515};
        10'd  436: lut_data <= {10'd15491};
        10'd  437: lut_data <= {10'd15468};
        10'd  438: lut_data <= {10'd15444};
        10'd  439: lut_data <= {10'd15420};
        10'd  440: lut_data <= {10'd15396};
        10'd  441: lut_data <= {10'd15371};
        10'd  442: lut_data <= {10'd15346};
        10'd  443: lut_data <= {10'd15321};
        10'd  444: lut_data <= {10'd15296};
        10'd  445: lut_data <= {10'd15270};
        10'd  446: lut_data <= {10'd15244};
        10'd  447: lut_data <= {10'd15218};
        10'd  448: lut_data <= {10'd15191};
        10'd  449: lut_data <= {10'd15164};
        10'd  450: lut_data <= {10'd15137};
        10'd  451: lut_data <= {10'd15109};
        10'd  452: lut_data <= {10'd15082};
        10'd  453: lut_data <= {10'd15053};
        10'd  454: lut_data <= {10'd15025};
        10'd  455: lut_data <= {10'd14996};
        10'd  456: lut_data <= {10'd14968};
        10'd  457: lut_data <= {10'd14938};
        10'd  458: lut_data <= {10'd14909};
        10'd  459: lut_data <= {10'd14879};
        10'd  460: lut_data <= {10'd14849};
        10'd  461: lut_data <= {10'd14819};
        10'd  462: lut_data <= {10'd14788};
        10'd  463: lut_data <= {10'd14757};
        10'd  464: lut_data <= {10'd14726};
        10'd  465: lut_data <= {10'd14694};
        10'd  466: lut_data <= {10'd14663};
        10'd  467: lut_data <= {10'd14631};
        10'd  468: lut_data <= {10'd14598};
        10'd  469: lut_data <= {10'd14566};
        10'd  470: lut_data <= {10'd14533};
        10'd  471: lut_data <= {10'd14500};
        10'd  472: lut_data <= {10'd14466};
        10'd  473: lut_data <= {10'd14433};
        10'd  474: lut_data <= {10'd14399};
        10'd  475: lut_data <= {10'd14364};
        10'd  476: lut_data <= {10'd14330};
        10'd  477: lut_data <= {10'd14295};
        10'd  478: lut_data <= {10'd14260};
        10'd  479: lut_data <= {10'd14225};
        10'd  480: lut_data <= {10'd14189};
        10'd  481: lut_data <= {10'd14153};
        10'd  482: lut_data <= {10'd14117};
        10'd  483: lut_data <= {10'd14081};
        10'd  484: lut_data <= {10'd14044};
        10'd  485: lut_data <= {10'd14007};
        10'd  486: lut_data <= {10'd13970};
        10'd  487: lut_data <= {10'd13932};
        10'd  488: lut_data <= {10'd13894};
        10'd  489: lut_data <= {10'd13856};
        10'd  490: lut_data <= {10'd13818};
        10'd  491: lut_data <= {10'd13780};
        10'd  492: lut_data <= {10'd13741};
        10'd  493: lut_data <= {10'd13702};
        10'd  494: lut_data <= {10'd13662};
        10'd  495: lut_data <= {10'd13623};
        10'd  496: lut_data <= {10'd13583};
        10'd  497: lut_data <= {10'd13543};
        10'd  498: lut_data <= {10'd13502};
        10'd  499: lut_data <= {10'd13462};
        10'd  500: lut_data <= {10'd13421};
        10'd  501: lut_data <= {10'd13380};
        10'd  502: lut_data <= {10'd13338};
        10'd  503: lut_data <= {10'd13297};
        10'd  504: lut_data <= {10'd13255};
        10'd  505: lut_data <= {10'd13213};
        10'd  506: lut_data <= {10'd13170};
        10'd  507: lut_data <= {10'd13128};
        10'd  508: lut_data <= {10'd13085};
        10'd  509: lut_data <= {10'd13042};
        10'd  510: lut_data <= {10'd12998};
        10'd  511: lut_data <= {10'd12955};
        10'd  512: lut_data <= {10'd12911};
        10'd  513: lut_data <= {10'd12867};
        10'd  514: lut_data <= {10'd12822};
        10'd  515: lut_data <= {10'd12778};
        10'd  516: lut_data <= {10'd12733};
        10'd  517: lut_data <= {10'd12688};
        10'd  518: lut_data <= {10'd12642};
        10'd  519: lut_data <= {10'd12597};
        10'd  520: lut_data <= {10'd12551};
        10'd  521: lut_data <= {10'd12505};
        10'd  522: lut_data <= {10'd12458};
        10'd  523: lut_data <= {10'd12412};
        10'd  524: lut_data <= {10'd12365};
        10'd  525: lut_data <= {10'd12318};
        10'd  526: lut_data <= {10'd12271};
        10'd  527: lut_data <= {10'd12223};
        10'd  528: lut_data <= {10'd12176};
        10'd  529: lut_data <= {10'd12128};
        10'd  530: lut_data <= {10'd12080};
        10'd  531: lut_data <= {10'd12031};
        10'd  532: lut_data <= {10'd11982};
        10'd  533: lut_data <= {10'd11934};
        10'd  534: lut_data <= {10'd11885};
        10'd  535: lut_data <= {10'd11835};
        10'd  536: lut_data <= {10'd11786};
        10'd  537: lut_data <= {10'd11736};
        10'd  538: lut_data <= {10'd11686};
        10'd  539: lut_data <= {10'd11636};
        10'd  540: lut_data <= {10'd11585};
        10'd  541: lut_data <= {10'd11535};
        10'd  542: lut_data <= {10'd11484};
        10'd  543: lut_data <= {10'd11433};
        10'd  544: lut_data <= {10'd11381};
        10'd  545: lut_data <= {10'd11330};
        10'd  546: lut_data <= {10'd11278};
        10'd  547: lut_data <= {10'd11226};
        10'd  548: lut_data <= {10'd11174};
        10'd  549: lut_data <= {10'd11121};
        10'd  550: lut_data <= {10'd11069};
        10'd  551: lut_data <= {10'd11016};
        10'd  552: lut_data <= {10'd10963};
        10'd  553: lut_data <= {10'd10910};
        10'd  554: lut_data <= {10'd10856};
        10'd  555: lut_data <= {10'd10803};
        10'd  556: lut_data <= {10'd10749};
        10'd  557: lut_data <= {10'd10695};
        10'd  558: lut_data <= {10'd10641};
        10'd  559: lut_data <= {10'd10586};
        10'd  560: lut_data <= {10'd10531};
        10'd  561: lut_data <= {10'd10477};
        10'd  562: lut_data <= {10'd10422};
        10'd  563: lut_data <= {10'd10366};
        10'd  564: lut_data <= {10'd10311};
        10'd  565: lut_data <= {10'd10255};
        10'd  566: lut_data <= {10'd10199};
        10'd  567: lut_data <= {10'd10143};
        10'd  568: lut_data <= {10'd10087};
        10'd  569: lut_data <= {10'd10031};
        10'd  570: lut_data <= {10'd09974};
        10'd  571: lut_data <= {10'd09917};
        10'd  572: lut_data <= {10'd09860};
        10'd  573: lut_data <= {10'd09803};
        10'd  574: lut_data <= {10'd09746};
        10'd  575: lut_data <= {10'd09688};
        10'd  576: lut_data <= {10'd09630};
        10'd  577: lut_data <= {10'd09572};
        10'd  578: lut_data <= {10'd09514};
        10'd  579: lut_data <= {10'd09456};
        10'd  580: lut_data <= {10'd09397};
        10'd  581: lut_data <= {10'd09339};
        10'd  582: lut_data <= {10'd09280};
        10'd  583: lut_data <= {10'd09221};
        10'd  584: lut_data <= {10'd09162};
        10'd  585: lut_data <= {10'd09102};
        10'd  586: lut_data <= {10'd09043};
        10'd  587: lut_data <= {10'd08983};
        10'd  588: lut_data <= {10'd08923};
        10'd  589: lut_data <= {10'd08863};
        10'd  590: lut_data <= {10'd08803};
        10'd  591: lut_data <= {10'd08743};
        10'd  592: lut_data <= {10'd08682};
        10'd  593: lut_data <= {10'd08621};
        10'd  594: lut_data <= {10'd08561};
        10'd  595: lut_data <= {10'd08500};
        10'd  596: lut_data <= {10'd08438};
        10'd  597: lut_data <= {10'd08377};
        10'd  598: lut_data <= {10'd08316};
        10'd  599: lut_data <= {10'd08254};
        10'd  600: lut_data <= {10'd08192};
        10'd  601: lut_data <= {10'd08130};
        10'd  602: lut_data <= {10'd08068};
        10'd  603: lut_data <= {10'd08006};
        10'd  604: lut_data <= {10'd07943};
        10'd  605: lut_data <= {10'd07881};
        10'd  606: lut_data <= {10'd07818};
        10'd  607: lut_data <= {10'd07755};
        10'd  608: lut_data <= {10'd07692};
        10'd  609: lut_data <= {10'd07629};
        10'd  610: lut_data <= {10'd07565};
        10'd  611: lut_data <= {10'd07502};
        10'd  612: lut_data <= {10'd07438};
        10'd  613: lut_data <= {10'd07374};
        10'd  614: lut_data <= {10'd07311};
        10'd  615: lut_data <= {10'd07246};
        10'd  616: lut_data <= {10'd07182};
        10'd  617: lut_data <= {10'd07118};
        10'd  618: lut_data <= {10'd07053};
        10'd  619: lut_data <= {10'd06989};
        10'd  620: lut_data <= {10'd06924};
        10'd  621: lut_data <= {10'd06859};
        10'd  622: lut_data <= {10'd06794};
        10'd  623: lut_data <= {10'd06729};
        10'd  624: lut_data <= {10'd06664};
        10'd  625: lut_data <= {10'd06599};
        10'd  626: lut_data <= {10'd06533};
        10'd  627: lut_data <= {10'd06467};
        10'd  628: lut_data <= {10'd06402};
        10'd  629: lut_data <= {10'd06336};
        10'd  630: lut_data <= {10'd06270};
        10'd  631: lut_data <= {10'd06204};
        10'd  632: lut_data <= {10'd06138};
        10'd  633: lut_data <= {10'd06071};
        10'd  634: lut_data <= {10'd06005};
        10'd  635: lut_data <= {10'd05938};
        10'd  636: lut_data <= {10'd05872};
        10'd  637: lut_data <= {10'd05805};
        10'd  638: lut_data <= {10'd05738};
        10'd  639: lut_data <= {10'd05671};
        10'd  640: lut_data <= {10'd05604};
        10'd  641: lut_data <= {10'd05536};
        10'd  642: lut_data <= {10'd05469};
        10'd  643: lut_data <= {10'd05402};
        10'd  644: lut_data <= {10'd05334};
        10'd  645: lut_data <= {10'd05266};
        10'd  646: lut_data <= {10'd05199};
        10'd  647: lut_data <= {10'd05131};
        10'd  648: lut_data <= {10'd05063};
        10'd  649: lut_data <= {10'd04995};
        10'd  650: lut_data <= {10'd04927};
        10'd  651: lut_data <= {10'd04859};
        10'd  652: lut_data <= {10'd04790};
        10'd  653: lut_data <= {10'd04722};
        10'd  654: lut_data <= {10'd04653};
        10'd  655: lut_data <= {10'd04585};
        10'd  656: lut_data <= {10'd04516};
        10'd  657: lut_data <= {10'd04447};
        10'd  658: lut_data <= {10'd04378};
        10'd  659: lut_data <= {10'd04310};
        10'd  660: lut_data <= {10'd04240};
        10'd  661: lut_data <= {10'd04171};
        10'd  662: lut_data <= {10'd04102};
        10'd  663: lut_data <= {10'd04033};
        10'd  664: lut_data <= {10'd03964};
        10'd  665: lut_data <= {10'd03894};
        10'd  666: lut_data <= {10'd03825};
        10'd  667: lut_data <= {10'd03755};
        10'd  668: lut_data <= {10'd03686};
        10'd  669: lut_data <= {10'd03616};
        10'd  670: lut_data <= {10'd03546};
        10'd  671: lut_data <= {10'd03476};
        10'd  672: lut_data <= {10'd03406};
        10'd  673: lut_data <= {10'd03336};
        10'd  674: lut_data <= {10'd03266};
        10'd  675: lut_data <= {10'd03196};
        10'd  676: lut_data <= {10'd03126};
        10'd  677: lut_data <= {10'd03056};
        10'd  678: lut_data <= {10'd02986};
        10'd  679: lut_data <= {10'd02915};
        10'd  680: lut_data <= {10'd02845};
        10'd  681: lut_data <= {10'd02775};
        10'd  682: lut_data <= {10'd02704};
        10'd  683: lut_data <= {10'd02634};
        10'd  684: lut_data <= {10'd02563};
        10'd  685: lut_data <= {10'd02492};
        10'd  686: lut_data <= {10'd02422};
        10'd  687: lut_data <= {10'd02351};
        10'd  688: lut_data <= {10'd02280};
        10'd  689: lut_data <= {10'd02209};
        10'd  690: lut_data <= {10'd02139};
        10'd  691: lut_data <= {10'd02068};
        10'd  692: lut_data <= {10'd01997};
        10'd  693: lut_data <= {10'd01926};
        10'd  694: lut_data <= {10'd01855};
        10'd  695: lut_data <= {10'd01784};
        10'd  696: lut_data <= {10'd01713};
        10'd  697: lut_data <= {10'd01641};
        10'd  698: lut_data <= {10'd01570};
        10'd  699: lut_data <= {10'd01499};
        10'd  700: lut_data <= {10'd01428};
        10'd  701: lut_data <= {10'd01357};
        10'd  702: lut_data <= {10'd01285};
        10'd  703: lut_data <= {10'd01214};
        10'd  704: lut_data <= {10'd01143};
        10'd  705: lut_data <= {10'd01072};
        10'd  706: lut_data <= {10'd01000};
        10'd  707: lut_data <= {10'd00929};
        10'd  708: lut_data <= {10'd00857};
        10'd  709: lut_data <= {10'd00786};
        10'd  710: lut_data <= {10'd00715};
        10'd  711: lut_data <= {10'd00643};
        10'd  712: lut_data <= {10'd00572};
        10'd  713: lut_data <= {10'd00500};
        10'd  714: lut_data <= {10'd00429};
        10'd  715: lut_data <= {10'd00357};
        10'd  716: lut_data <= {10'd00286};
        10'd  717: lut_data <= {10'd00214};
        10'd  718: lut_data <= {10'd00143};
        10'd  719: lut_data <= {10'd00071};
        10'd  720: lut_data <= {10'd00000};
        10'd  721: lut_data <= {-10'd00071};
        10'd  722: lut_data <= {-10'd00143};
        10'd  723: lut_data <= {-10'd00214};
        10'd  724: lut_data <= {-10'd00286};
        10'd  725: lut_data <= {-10'd00357};
        10'd  726: lut_data <= {-10'd00429};
        10'd  727: lut_data <= {-10'd00500};
        10'd  728: lut_data <= {-10'd00572};
        10'd  729: lut_data <= {-10'd00643};
        10'd  730: lut_data <= {-10'd00715};
        10'd  731: lut_data <= {-10'd00786};
        10'd  732: lut_data <= {-10'd00857};
        10'd  733: lut_data <= {-10'd00929};
        10'd  734: lut_data <= {-10'd01000};
        10'd  735: lut_data <= {-10'd01072};
        10'd  736: lut_data <= {-10'd01143};
        10'd  737: lut_data <= {-10'd01214};
        10'd  738: lut_data <= {-10'd01285};
        10'd  739: lut_data <= {-10'd01357};
        10'd  740: lut_data <= {-10'd01428};
        10'd  741: lut_data <= {-10'd01499};
        10'd  742: lut_data <= {-10'd01570};
        10'd  743: lut_data <= {-10'd01641};
        10'd  744: lut_data <= {-10'd01713};
        10'd  745: lut_data <= {-10'd01784};
        10'd  746: lut_data <= {-10'd01855};
        10'd  747: lut_data <= {-10'd01926};
        10'd  748: lut_data <= {-10'd01997};
        10'd  749: lut_data <= {-10'd02068};
        10'd  750: lut_data <= {-10'd02139};
        10'd  751: lut_data <= {-10'd02209};
        10'd  752: lut_data <= {-10'd02280};
        10'd  753: lut_data <= {-10'd02351};
        10'd  754: lut_data <= {-10'd02422};
        10'd  755: lut_data <= {-10'd02492};
        10'd  756: lut_data <= {-10'd02563};
        10'd  757: lut_data <= {-10'd02634};
        10'd  758: lut_data <= {-10'd02704};
        10'd  759: lut_data <= {-10'd02775};
        10'd  760: lut_data <= {-10'd02845};
        10'd  761: lut_data <= {-10'd02915};
        10'd  762: lut_data <= {-10'd02986};
        10'd  763: lut_data <= {-10'd03056};
        10'd  764: lut_data <= {-10'd03126};
        10'd  765: lut_data <= {-10'd03196};
        10'd  766: lut_data <= {-10'd03266};
        10'd  767: lut_data <= {-10'd03336};
        10'd  768: lut_data <= {-10'd03406};
        10'd  769: lut_data <= {-10'd03476};
        10'd  770: lut_data <= {-10'd03546};
        10'd  771: lut_data <= {-10'd03616};
        10'd  772: lut_data <= {-10'd03686};
        10'd  773: lut_data <= {-10'd03755};
        10'd  774: lut_data <= {-10'd03825};
        10'd  775: lut_data <= {-10'd03894};
        10'd  776: lut_data <= {-10'd03964};
        10'd  777: lut_data <= {-10'd04033};
        10'd  778: lut_data <= {-10'd04102};
        10'd  779: lut_data <= {-10'd04171};
        10'd  780: lut_data <= {-10'd04240};
        10'd  781: lut_data <= {-10'd04310};
        10'd  782: lut_data <= {-10'd04378};
        10'd  783: lut_data <= {-10'd04447};
        10'd  784: lut_data <= {-10'd04516};
        10'd  785: lut_data <= {-10'd04585};
        10'd  786: lut_data <= {-10'd04653};
        10'd  787: lut_data <= {-10'd04722};
        10'd  788: lut_data <= {-10'd04790};
        10'd  789: lut_data <= {-10'd04859};
        10'd  790: lut_data <= {-10'd04927};
        10'd  791: lut_data <= {-10'd04995};
        10'd  792: lut_data <= {-10'd05063};
        10'd  793: lut_data <= {-10'd05131};
        10'd  794: lut_data <= {-10'd05199};
        10'd  795: lut_data <= {-10'd05266};
        10'd  796: lut_data <= {-10'd05334};
        10'd  797: lut_data <= {-10'd05402};
        10'd  798: lut_data <= {-10'd05469};
        10'd  799: lut_data <= {-10'd05536};
        10'd  800: lut_data <= {-10'd05604};
        10'd  801: lut_data <= {-10'd05671};
        10'd  802: lut_data <= {-10'd05738};
        10'd  803: lut_data <= {-10'd05805};
        10'd  804: lut_data <= {-10'd05872};
        10'd  805: lut_data <= {-10'd05938};
        10'd  806: lut_data <= {-10'd06005};
        10'd  807: lut_data <= {-10'd06071};
        10'd  808: lut_data <= {-10'd06138};
        10'd  809: lut_data <= {-10'd06204};
        10'd  810: lut_data <= {-10'd06270};
        10'd  811: lut_data <= {-10'd06336};
        10'd  812: lut_data <= {-10'd06402};
        10'd  813: lut_data <= {-10'd06467};
        10'd  814: lut_data <= {-10'd06533};
        10'd  815: lut_data <= {-10'd06599};
        10'd  816: lut_data <= {-10'd06664};
        10'd  817: lut_data <= {-10'd06729};
        10'd  818: lut_data <= {-10'd06794};
        10'd  819: lut_data <= {-10'd06859};
        10'd  820: lut_data <= {-10'd06924};
        10'd  821: lut_data <= {-10'd06989};
        10'd  822: lut_data <= {-10'd07053};
        10'd  823: lut_data <= {-10'd07118};
        10'd  824: lut_data <= {-10'd07182};
        10'd  825: lut_data <= {-10'd07246};
        10'd  826: lut_data <= {-10'd07311};
        10'd  827: lut_data <= {-10'd07374};
        10'd  828: lut_data <= {-10'd07438};
        10'd  829: lut_data <= {-10'd07502};
        10'd  830: lut_data <= {-10'd07565};
        10'd  831: lut_data <= {-10'd07629};
        10'd  832: lut_data <= {-10'd07692};
        10'd  833: lut_data <= {-10'd07755};
        10'd  834: lut_data <= {-10'd07818};
        10'd  835: lut_data <= {-10'd07881};
        10'd  836: lut_data <= {-10'd07943};
        10'd  837: lut_data <= {-10'd08006};
        10'd  838: lut_data <= {-10'd08068};
        10'd  839: lut_data <= {-10'd08130};
        10'd  840: lut_data <= {-10'd08192};
        10'd  841: lut_data <= {-10'd08254};
        10'd  842: lut_data <= {-10'd08316};
        10'd  843: lut_data <= {-10'd08377};
        10'd  844: lut_data <= {-10'd08438};
        10'd  845: lut_data <= {-10'd08500};
        10'd  846: lut_data <= {-10'd08561};
        10'd  847: lut_data <= {-10'd08621};
        10'd  848: lut_data <= {-10'd08682};
        10'd  849: lut_data <= {-10'd08743};
        10'd  850: lut_data <= {-10'd08803};
        10'd  851: lut_data <= {-10'd08863};
        10'd  852: lut_data <= {-10'd08923};
        10'd  853: lut_data <= {-10'd08983};
        10'd  854: lut_data <= {-10'd09043};
        10'd  855: lut_data <= {-10'd09102};
        10'd  856: lut_data <= {-10'd09162};
        10'd  857: lut_data <= {-10'd09221};
        10'd  858: lut_data <= {-10'd09280};
        10'd  859: lut_data <= {-10'd09339};
        10'd  860: lut_data <= {-10'd09397};
        10'd  861: lut_data <= {-10'd09456};
        10'd  862: lut_data <= {-10'd09514};
        10'd  863: lut_data <= {-10'd09572};
        10'd  864: lut_data <= {-10'd09630};
        10'd  865: lut_data <= {-10'd09688};
        10'd  866: lut_data <= {-10'd09746};
        10'd  867: lut_data <= {-10'd09803};
        10'd  868: lut_data <= {-10'd09860};
        10'd  869: lut_data <= {-10'd09917};
        10'd  870: lut_data <= {-10'd09974};
        10'd  871: lut_data <= {-10'd10031};
        10'd  872: lut_data <= {-10'd10087};
        10'd  873: lut_data <= {-10'd10143};
        10'd  874: lut_data <= {-10'd10199};
        10'd  875: lut_data <= {-10'd10255};
        10'd  876: lut_data <= {-10'd10311};
        10'd  877: lut_data <= {-10'd10366};
        10'd  878: lut_data <= {-10'd10422};
        10'd  879: lut_data <= {-10'd10477};
        10'd  880: lut_data <= {-10'd10531};
        10'd  881: lut_data <= {-10'd10586};
        10'd  882: lut_data <= {-10'd10641};
        10'd  883: lut_data <= {-10'd10695};
        10'd  884: lut_data <= {-10'd10749};
        10'd  885: lut_data <= {-10'd10803};
        10'd  886: lut_data <= {-10'd10856};
        10'd  887: lut_data <= {-10'd10910};
        10'd  888: lut_data <= {-10'd10963};
        10'd  889: lut_data <= {-10'd11016};
        10'd  890: lut_data <= {-10'd11069};
        10'd  891: lut_data <= {-10'd11121};
        10'd  892: lut_data <= {-10'd11174};
        10'd  893: lut_data <= {-10'd11226};
        10'd  894: lut_data <= {-10'd11278};
        10'd  895: lut_data <= {-10'd11330};
        10'd  896: lut_data <= {-10'd11381};
        10'd  897: lut_data <= {-10'd11433};
        10'd  898: lut_data <= {-10'd11484};
        10'd  899: lut_data <= {-10'd11535};
        10'd  900: lut_data <= {-10'd11585};
        10'd  901: lut_data <= {-10'd11636};
        10'd  902: lut_data <= {-10'd11686};
        10'd  903: lut_data <= {-10'd11736};
        10'd  904: lut_data <= {-10'd11786};
        10'd  905: lut_data <= {-10'd11835};
        10'd  906: lut_data <= {-10'd11885};
        10'd  907: lut_data <= {-10'd11934};
        10'd  908: lut_data <= {-10'd11982};
        10'd  909: lut_data <= {-10'd12031};
        10'd  910: lut_data <= {-10'd12080};
        10'd  911: lut_data <= {-10'd12128};
        10'd  912: lut_data <= {-10'd12176};
        10'd  913: lut_data <= {-10'd12223};
        10'd  914: lut_data <= {-10'd12271};
        10'd  915: lut_data <= {-10'd12318};
        10'd  916: lut_data <= {-10'd12365};
        10'd  917: lut_data <= {-10'd12412};
        10'd  918: lut_data <= {-10'd12458};
        10'd  919: lut_data <= {-10'd12505};
        10'd  920: lut_data <= {-10'd12551};
        10'd  921: lut_data <= {-10'd12597};
        10'd  922: lut_data <= {-10'd12642};
        10'd  923: lut_data <= {-10'd12688};
        10'd  924: lut_data <= {-10'd12733};
        10'd  925: lut_data <= {-10'd12778};
        10'd  926: lut_data <= {-10'd12822};
        10'd  927: lut_data <= {-10'd12867};
        10'd  928: lut_data <= {-10'd12911};
        10'd  929: lut_data <= {-10'd12955};
        10'd  930: lut_data <= {-10'd12998};
        10'd  931: lut_data <= {-10'd13042};
        10'd  932: lut_data <= {-10'd13085};
        10'd  933: lut_data <= {-10'd13128};
        10'd  934: lut_data <= {-10'd13170};
        10'd  935: lut_data <= {-10'd13213};
        10'd  936: lut_data <= {-10'd13255};
        10'd  937: lut_data <= {-10'd13297};
        10'd  938: lut_data <= {-10'd13338};
        10'd  939: lut_data <= {-10'd13380};
        10'd  940: lut_data <= {-10'd13421};
        10'd  941: lut_data <= {-10'd13462};
        10'd  942: lut_data <= {-10'd13502};
        10'd  943: lut_data <= {-10'd13543};
        10'd  944: lut_data <= {-10'd13583};
        10'd  945: lut_data <= {-10'd13623};
        10'd  946: lut_data <= {-10'd13662};
        10'd  947: lut_data <= {-10'd13702};
        10'd  948: lut_data <= {-10'd13741};
        10'd  949: lut_data <= {-10'd13780};
        10'd  950: lut_data <= {-10'd13818};
        10'd  951: lut_data <= {-10'd13856};
        10'd  952: lut_data <= {-10'd13894};
        10'd  953: lut_data <= {-10'd13932};
        10'd  954: lut_data <= {-10'd13970};
        10'd  955: lut_data <= {-10'd14007};
        10'd  956: lut_data <= {-10'd14044};
        10'd  957: lut_data <= {-10'd14081};
        10'd  958: lut_data <= {-10'd14117};
        10'd  959: lut_data <= {-10'd14153};
        10'd  960: lut_data <= {-10'd14189};
        10'd  961: lut_data <= {-10'd14225};
        10'd  962: lut_data <= {-10'd14260};
        10'd  963: lut_data <= {-10'd14295};
        10'd  964: lut_data <= {-10'd14330};
        10'd  965: lut_data <= {-10'd14364};
        10'd  966: lut_data <= {-10'd14399};
        10'd  967: lut_data <= {-10'd14433};
        10'd  968: lut_data <= {-10'd14466};
        10'd  969: lut_data <= {-10'd14500};
        10'd  970: lut_data <= {-10'd14533};
        10'd  971: lut_data <= {-10'd14566};
        10'd  972: lut_data <= {-10'd14598};
        10'd  973: lut_data <= {-10'd14631};
        10'd  974: lut_data <= {-10'd14663};
        10'd  975: lut_data <= {-10'd14694};
        10'd  976: lut_data <= {-10'd14726};
        10'd  977: lut_data <= {-10'd14757};
        10'd  978: lut_data <= {-10'd14788};
        10'd  979: lut_data <= {-10'd14819};
        10'd  980: lut_data <= {-10'd14849};
        10'd  981: lut_data <= {-10'd14879};
        10'd  982: lut_data <= {-10'd14909};
        10'd  983: lut_data <= {-10'd14938};
        10'd  984: lut_data <= {-10'd14968};
        10'd  985: lut_data <= {-10'd14996};
        10'd  986: lut_data <= {-10'd15025};
        10'd  987: lut_data <= {-10'd15053};
        10'd  988: lut_data <= {-10'd15082};
        10'd  989: lut_data <= {-10'd15109};
        10'd  990: lut_data <= {-10'd15137};
        10'd  991: lut_data <= {-10'd15164};
        10'd  992: lut_data <= {-10'd15191};
        10'd  993: lut_data <= {-10'd15218};
        10'd  994: lut_data <= {-10'd15244};
        10'd  995: lut_data <= {-10'd15270};
        10'd  996: lut_data <= {-10'd15296};
        10'd  997: lut_data <= {-10'd15321};
        10'd  998: lut_data <= {-10'd15346};
        10'd  999: lut_data <= {-10'd15371};
        10'd 1000: lut_data <= {-10'd15396};
        10'd 1001: lut_data <= {-10'd15420};
        10'd 1002: lut_data <= {-10'd15444};
        10'd 1003: lut_data <= {-10'd15468};
        10'd 1004: lut_data <= {-10'd15491};
        10'd 1005: lut_data <= {-10'd15515};
        10'd 1006: lut_data <= {-10'd15537};
        10'd 1007: lut_data <= {-10'd15560};
        10'd 1008: lut_data <= {-10'd15582};
        10'd 1009: lut_data <= {-10'd15604};
        10'd 1010: lut_data <= {-10'd15626};
        10'd 1011: lut_data <= {-10'd15647};
        10'd 1012: lut_data <= {-10'd15668};
        10'd 1013: lut_data <= {-10'd15689};
        10'd 1014: lut_data <= {-10'd15709};
        10'd 1015: lut_data <= {-10'd15729};
        10'd 1016: lut_data <= {-10'd15749};
        10'd 1017: lut_data <= {-10'd15769};
        10'd 1018: lut_data <= {-10'd15788};
        10'd 1019: lut_data <= {-10'd15807};
        10'd 1020: lut_data <= {-10'd15826};
        10'd 1021: lut_data <= {-10'd15844};
        10'd 1022: lut_data <= {-10'd15862};
        10'd 1023: lut_data <= {-10'd15880};
        10'd 1024: lut_data <= {-10'd15897};
        10'd 1025: lut_data <= {-10'd15914};
        10'd 1026: lut_data <= {-10'd15931};
        10'd 1027: lut_data <= {-10'd15948};
        10'd 1028: lut_data <= {-10'd15964};
        10'd 1029: lut_data <= {-10'd15980};
        10'd 1030: lut_data <= {-10'd15996};
        10'd 1031: lut_data <= {-10'd16011};
        10'd 1032: lut_data <= {-10'd16026};
        10'd 1033: lut_data <= {-10'd16041};
        10'd 1034: lut_data <= {-10'd16055};
        10'd 1035: lut_data <= {-10'd16069};
        10'd 1036: lut_data <= {-10'd16083};
        10'd 1037: lut_data <= {-10'd16096};
        10'd 1038: lut_data <= {-10'd16110};
        10'd 1039: lut_data <= {-10'd16123};
        10'd 1040: lut_data <= {-10'd16135};
        10'd 1041: lut_data <= {-10'd16147};
        10'd 1042: lut_data <= {-10'd16159};
        10'd 1043: lut_data <= {-10'd16171};
        10'd 1044: lut_data <= {-10'd16182};
        10'd 1045: lut_data <= {-10'd16193};
        10'd 1046: lut_data <= {-10'd16204};
        10'd 1047: lut_data <= {-10'd16214};
        10'd 1048: lut_data <= {-10'd16225};
        10'd 1049: lut_data <= {-10'd16234};
        10'd 1050: lut_data <= {-10'd16244};
        10'd 1051: lut_data <= {-10'd16253};
        10'd 1052: lut_data <= {-10'd16262};
        10'd 1053: lut_data <= {-10'd16270};
        10'd 1054: lut_data <= {-10'd16279};
        10'd 1055: lut_data <= {-10'd16287};
        10'd 1056: lut_data <= {-10'd16294};
        10'd 1057: lut_data <= {-10'd16302};
        10'd 1058: lut_data <= {-10'd16309};
        10'd 1059: lut_data <= {-10'd16315};
        10'd 1060: lut_data <= {-10'd16322};
        10'd 1061: lut_data <= {-10'd16328};
        10'd 1062: lut_data <= {-10'd16333};
        10'd 1063: lut_data <= {-10'd16339};
        10'd 1064: lut_data <= {-10'd16344};
        10'd 1065: lut_data <= {-10'd16349};
        10'd 1066: lut_data <= {-10'd16353};
        10'd 1067: lut_data <= {-10'd16358};
        10'd 1068: lut_data <= {-10'd16362};
        10'd 1069: lut_data <= {-10'd16365};
        10'd 1070: lut_data <= {-10'd16368};
        10'd 1071: lut_data <= {-10'd16371};
        10'd 1072: lut_data <= {-10'd16374};
        10'd 1073: lut_data <= {-10'd16376};
        10'd 1074: lut_data <= {-10'd16378};
        10'd 1075: lut_data <= {-10'd16380};
        10'd 1076: lut_data <= {-10'd16382};
        10'd 1077: lut_data <= {-10'd16383};
        10'd 1078: lut_data <= {-10'd16383};
        10'd 1079: lut_data <= {-10'd16384};
        10'd 1080: lut_data <= {-10'd16384};
        10'd 1081: lut_data <= {-10'd16384};
        10'd 1082: lut_data <= {-10'd16383};
        10'd 1083: lut_data <= {-10'd16383};
        10'd 1084: lut_data <= {-10'd16382};
        10'd 1085: lut_data <= {-10'd16380};
        10'd 1086: lut_data <= {-10'd16378};
        10'd 1087: lut_data <= {-10'd16376};
        10'd 1088: lut_data <= {-10'd16374};
        10'd 1089: lut_data <= {-10'd16371};
        10'd 1090: lut_data <= {-10'd16368};
        10'd 1091: lut_data <= {-10'd16365};
        10'd 1092: lut_data <= {-10'd16362};
        10'd 1093: lut_data <= {-10'd16358};
        10'd 1094: lut_data <= {-10'd16353};
        10'd 1095: lut_data <= {-10'd16349};
        10'd 1096: lut_data <= {-10'd16344};
        10'd 1097: lut_data <= {-10'd16339};
        10'd 1098: lut_data <= {-10'd16333};
        10'd 1099: lut_data <= {-10'd16328};
        10'd 1100: lut_data <= {-10'd16322};
        10'd 1101: lut_data <= {-10'd16315};
        10'd 1102: lut_data <= {-10'd16309};
        10'd 1103: lut_data <= {-10'd16302};
        10'd 1104: lut_data <= {-10'd16294};
        10'd 1105: lut_data <= {-10'd16287};
        10'd 1106: lut_data <= {-10'd16279};
        10'd 1107: lut_data <= {-10'd16270};
        10'd 1108: lut_data <= {-10'd16262};
        10'd 1109: lut_data <= {-10'd16253};
        10'd 1110: lut_data <= {-10'd16244};
        10'd 1111: lut_data <= {-10'd16234};
        10'd 1112: lut_data <= {-10'd16225};
        10'd 1113: lut_data <= {-10'd16214};
        10'd 1114: lut_data <= {-10'd16204};
        10'd 1115: lut_data <= {-10'd16193};
        10'd 1116: lut_data <= {-10'd16182};
        10'd 1117: lut_data <= {-10'd16171};
        10'd 1118: lut_data <= {-10'd16159};
        10'd 1119: lut_data <= {-10'd16147};
        10'd 1120: lut_data <= {-10'd16135};
        10'd 1121: lut_data <= {-10'd16123};
        10'd 1122: lut_data <= {-10'd16110};
        10'd 1123: lut_data <= {-10'd16096};
        10'd 1124: lut_data <= {-10'd16083};
        10'd 1125: lut_data <= {-10'd16069};
        10'd 1126: lut_data <= {-10'd16055};
        10'd 1127: lut_data <= {-10'd16041};
        10'd 1128: lut_data <= {-10'd16026};
        10'd 1129: lut_data <= {-10'd16011};
        10'd 1130: lut_data <= {-10'd15996};
        10'd 1131: lut_data <= {-10'd15980};
        10'd 1132: lut_data <= {-10'd15964};
        10'd 1133: lut_data <= {-10'd15948};
        10'd 1134: lut_data <= {-10'd15931};
        10'd 1135: lut_data <= {-10'd15914};
        10'd 1136: lut_data <= {-10'd15897};
        10'd 1137: lut_data <= {-10'd15880};
        10'd 1138: lut_data <= {-10'd15862};
        10'd 1139: lut_data <= {-10'd15844};
        10'd 1140: lut_data <= {-10'd15826};
        10'd 1141: lut_data <= {-10'd15807};
        10'd 1142: lut_data <= {-10'd15788};
        10'd 1143: lut_data <= {-10'd15769};
        10'd 1144: lut_data <= {-10'd15749};
        10'd 1145: lut_data <= {-10'd15729};
        10'd 1146: lut_data <= {-10'd15709};
        10'd 1147: lut_data <= {-10'd15689};
        10'd 1148: lut_data <= {-10'd15668};
        10'd 1149: lut_data <= {-10'd15647};
        10'd 1150: lut_data <= {-10'd15626};
        10'd 1151: lut_data <= {-10'd15604};
        10'd 1152: lut_data <= {-10'd15582};
        10'd 1153: lut_data <= {-10'd15560};
        10'd 1154: lut_data <= {-10'd15537};
        10'd 1155: lut_data <= {-10'd15515};
        10'd 1156: lut_data <= {-10'd15491};
        10'd 1157: lut_data <= {-10'd15468};
        10'd 1158: lut_data <= {-10'd15444};
        10'd 1159: lut_data <= {-10'd15420};
        10'd 1160: lut_data <= {-10'd15396};
        10'd 1161: lut_data <= {-10'd15371};
        10'd 1162: lut_data <= {-10'd15346};
        10'd 1163: lut_data <= {-10'd15321};
        10'd 1164: lut_data <= {-10'd15296};
        10'd 1165: lut_data <= {-10'd15270};
        10'd 1166: lut_data <= {-10'd15244};
        10'd 1167: lut_data <= {-10'd15218};
        10'd 1168: lut_data <= {-10'd15191};
        10'd 1169: lut_data <= {-10'd15164};
        10'd 1170: lut_data <= {-10'd15137};
        10'd 1171: lut_data <= {-10'd15109};
        10'd 1172: lut_data <= {-10'd15082};
        10'd 1173: lut_data <= {-10'd15053};
        10'd 1174: lut_data <= {-10'd15025};
        10'd 1175: lut_data <= {-10'd14996};
        10'd 1176: lut_data <= {-10'd14968};
        10'd 1177: lut_data <= {-10'd14938};
        10'd 1178: lut_data <= {-10'd14909};
        10'd 1179: lut_data <= {-10'd14879};
        10'd 1180: lut_data <= {-10'd14849};
        10'd 1181: lut_data <= {-10'd14819};
        10'd 1182: lut_data <= {-10'd14788};
        10'd 1183: lut_data <= {-10'd14757};
        10'd 1184: lut_data <= {-10'd14726};
        10'd 1185: lut_data <= {-10'd14694};
        10'd 1186: lut_data <= {-10'd14663};
        10'd 1187: lut_data <= {-10'd14631};
        10'd 1188: lut_data <= {-10'd14598};
        10'd 1189: lut_data <= {-10'd14566};
        10'd 1190: lut_data <= {-10'd14533};
        10'd 1191: lut_data <= {-10'd14500};
        10'd 1192: lut_data <= {-10'd14466};
        10'd 1193: lut_data <= {-10'd14433};
        10'd 1194: lut_data <= {-10'd14399};
        10'd 1195: lut_data <= {-10'd14364};
        10'd 1196: lut_data <= {-10'd14330};
        10'd 1197: lut_data <= {-10'd14295};
        10'd 1198: lut_data <= {-10'd14260};
        10'd 1199: lut_data <= {-10'd14225};
        10'd 1200: lut_data <= {-10'd14189};
        10'd 1201: lut_data <= {-10'd14153};
        10'd 1202: lut_data <= {-10'd14117};
        10'd 1203: lut_data <= {-10'd14081};
        10'd 1204: lut_data <= {-10'd14044};
        10'd 1205: lut_data <= {-10'd14007};
        10'd 1206: lut_data <= {-10'd13970};
        10'd 1207: lut_data <= {-10'd13932};
        10'd 1208: lut_data <= {-10'd13894};
        10'd 1209: lut_data <= {-10'd13856};
        10'd 1210: lut_data <= {-10'd13818};
        10'd 1211: lut_data <= {-10'd13780};
        10'd 1212: lut_data <= {-10'd13741};
        10'd 1213: lut_data <= {-10'd13702};
        10'd 1214: lut_data <= {-10'd13662};
        10'd 1215: lut_data <= {-10'd13623};
        10'd 1216: lut_data <= {-10'd13583};
        10'd 1217: lut_data <= {-10'd13543};
        10'd 1218: lut_data <= {-10'd13502};
        10'd 1219: lut_data <= {-10'd13462};
        10'd 1220: lut_data <= {-10'd13421};
        10'd 1221: lut_data <= {-10'd13380};
        10'd 1222: lut_data <= {-10'd13338};
        10'd 1223: lut_data <= {-10'd13297};
        10'd 1224: lut_data <= {-10'd13255};
        10'd 1225: lut_data <= {-10'd13213};
        10'd 1226: lut_data <= {-10'd13170};
        10'd 1227: lut_data <= {-10'd13128};
        10'd 1228: lut_data <= {-10'd13085};
        10'd 1229: lut_data <= {-10'd13042};
        10'd 1230: lut_data <= {-10'd12998};
        10'd 1231: lut_data <= {-10'd12955};
        10'd 1232: lut_data <= {-10'd12911};
        10'd 1233: lut_data <= {-10'd12867};
        10'd 1234: lut_data <= {-10'd12822};
        10'd 1235: lut_data <= {-10'd12778};
        10'd 1236: lut_data <= {-10'd12733};
        10'd 1237: lut_data <= {-10'd12688};
        10'd 1238: lut_data <= {-10'd12642};
        10'd 1239: lut_data <= {-10'd12597};
        10'd 1240: lut_data <= {-10'd12551};
        10'd 1241: lut_data <= {-10'd12505};
        10'd 1242: lut_data <= {-10'd12458};
        10'd 1243: lut_data <= {-10'd12412};
        10'd 1244: lut_data <= {-10'd12365};
        10'd 1245: lut_data <= {-10'd12318};
        10'd 1246: lut_data <= {-10'd12271};
        10'd 1247: lut_data <= {-10'd12223};
        10'd 1248: lut_data <= {-10'd12176};
        10'd 1249: lut_data <= {-10'd12128};
        10'd 1250: lut_data <= {-10'd12080};
        10'd 1251: lut_data <= {-10'd12031};
        10'd 1252: lut_data <= {-10'd11982};
        10'd 1253: lut_data <= {-10'd11934};
        10'd 1254: lut_data <= {-10'd11885};
        10'd 1255: lut_data <= {-10'd11835};
        10'd 1256: lut_data <= {-10'd11786};
        10'd 1257: lut_data <= {-10'd11736};
        10'd 1258: lut_data <= {-10'd11686};
        10'd 1259: lut_data <= {-10'd11636};
        10'd 1260: lut_data <= {-10'd11585};
        10'd 1261: lut_data <= {-10'd11535};
        10'd 1262: lut_data <= {-10'd11484};
        10'd 1263: lut_data <= {-10'd11433};
        10'd 1264: lut_data <= {-10'd11381};
        10'd 1265: lut_data <= {-10'd11330};
        10'd 1266: lut_data <= {-10'd11278};
        10'd 1267: lut_data <= {-10'd11226};
        10'd 1268: lut_data <= {-10'd11174};
        10'd 1269: lut_data <= {-10'd11121};
        10'd 1270: lut_data <= {-10'd11069};
        10'd 1271: lut_data <= {-10'd11016};
        10'd 1272: lut_data <= {-10'd10963};
        10'd 1273: lut_data <= {-10'd10910};
        10'd 1274: lut_data <= {-10'd10856};
        10'd 1275: lut_data <= {-10'd10803};
        10'd 1276: lut_data <= {-10'd10749};
        10'd 1277: lut_data <= {-10'd10695};
        10'd 1278: lut_data <= {-10'd10641};
        10'd 1279: lut_data <= {-10'd10586};
        10'd 1280: lut_data <= {-10'd10531};
        10'd 1281: lut_data <= {-10'd10477};
        10'd 1282: lut_data <= {-10'd10422};
        10'd 1283: lut_data <= {-10'd10366};
        10'd 1284: lut_data <= {-10'd10311};
        10'd 1285: lut_data <= {-10'd10255};
        10'd 1286: lut_data <= {-10'd10199};
        10'd 1287: lut_data <= {-10'd10143};
        10'd 1288: lut_data <= {-10'd10087};
        10'd 1289: lut_data <= {-10'd10031};
        10'd 1290: lut_data <= {-10'd09974};
        10'd 1291: lut_data <= {-10'd09917};
        10'd 1292: lut_data <= {-10'd09860};
        10'd 1293: lut_data <= {-10'd09803};
        10'd 1294: lut_data <= {-10'd09746};
        10'd 1295: lut_data <= {-10'd09688};
        10'd 1296: lut_data <= {-10'd09630};
        10'd 1297: lut_data <= {-10'd09572};
        10'd 1298: lut_data <= {-10'd09514};
        10'd 1299: lut_data <= {-10'd09456};
        10'd 1300: lut_data <= {-10'd09397};
        10'd 1301: lut_data <= {-10'd09339};
        10'd 1302: lut_data <= {-10'd09280};
        10'd 1303: lut_data <= {-10'd09221};
        10'd 1304: lut_data <= {-10'd09162};
        10'd 1305: lut_data <= {-10'd09102};
        10'd 1306: lut_data <= {-10'd09043};
        10'd 1307: lut_data <= {-10'd08983};
        10'd 1308: lut_data <= {-10'd08923};
        10'd 1309: lut_data <= {-10'd08863};
        10'd 1310: lut_data <= {-10'd08803};
        10'd 1311: lut_data <= {-10'd08743};
        10'd 1312: lut_data <= {-10'd08682};
        10'd 1313: lut_data <= {-10'd08621};
        10'd 1314: lut_data <= {-10'd08561};
        10'd 1315: lut_data <= {-10'd08500};
        10'd 1316: lut_data <= {-10'd08438};
        10'd 1317: lut_data <= {-10'd08377};
        10'd 1318: lut_data <= {-10'd08316};
        10'd 1319: lut_data <= {-10'd08254};
        10'd 1320: lut_data <= {-10'd08192};
        10'd 1321: lut_data <= {-10'd08130};
        10'd 1322: lut_data <= {-10'd08068};
        10'd 1323: lut_data <= {-10'd08006};
        10'd 1324: lut_data <= {-10'd07943};
        10'd 1325: lut_data <= {-10'd07881};
        10'd 1326: lut_data <= {-10'd07818};
        10'd 1327: lut_data <= {-10'd07755};
        10'd 1328: lut_data <= {-10'd07692};
        10'd 1329: lut_data <= {-10'd07629};
        10'd 1330: lut_data <= {-10'd07565};
        10'd 1331: lut_data <= {-10'd07502};
        10'd 1332: lut_data <= {-10'd07438};
        10'd 1333: lut_data <= {-10'd07374};
        10'd 1334: lut_data <= {-10'd07311};
        10'd 1335: lut_data <= {-10'd07246};
        10'd 1336: lut_data <= {-10'd07182};
        10'd 1337: lut_data <= {-10'd07118};
        10'd 1338: lut_data <= {-10'd07053};
        10'd 1339: lut_data <= {-10'd06989};
        10'd 1340: lut_data <= {-10'd06924};
        10'd 1341: lut_data <= {-10'd06859};
        10'd 1342: lut_data <= {-10'd06794};
        10'd 1343: lut_data <= {-10'd06729};
        10'd 1344: lut_data <= {-10'd06664};
        10'd 1345: lut_data <= {-10'd06599};
        10'd 1346: lut_data <= {-10'd06533};
        10'd 1347: lut_data <= {-10'd06467};
        10'd 1348: lut_data <= {-10'd06402};
        10'd 1349: lut_data <= {-10'd06336};
        10'd 1350: lut_data <= {-10'd06270};
        10'd 1351: lut_data <= {-10'd06204};
        10'd 1352: lut_data <= {-10'd06138};
        10'd 1353: lut_data <= {-10'd06071};
        10'd 1354: lut_data <= {-10'd06005};
        10'd 1355: lut_data <= {-10'd05938};
        10'd 1356: lut_data <= {-10'd05872};
        10'd 1357: lut_data <= {-10'd05805};
        10'd 1358: lut_data <= {-10'd05738};
        10'd 1359: lut_data <= {-10'd05671};
        10'd 1360: lut_data <= {-10'd05604};
        10'd 1361: lut_data <= {-10'd05536};
        10'd 1362: lut_data <= {-10'd05469};
        10'd 1363: lut_data <= {-10'd05402};
        10'd 1364: lut_data <= {-10'd05334};
        10'd 1365: lut_data <= {-10'd05266};
        10'd 1366: lut_data <= {-10'd05199};
        10'd 1367: lut_data <= {-10'd05131};
        10'd 1368: lut_data <= {-10'd05063};
        10'd 1369: lut_data <= {-10'd04995};
        10'd 1370: lut_data <= {-10'd04927};
        10'd 1371: lut_data <= {-10'd04859};
        10'd 1372: lut_data <= {-10'd04790};
        10'd 1373: lut_data <= {-10'd04722};
        10'd 1374: lut_data <= {-10'd04653};
        10'd 1375: lut_data <= {-10'd04585};
        10'd 1376: lut_data <= {-10'd04516};
        10'd 1377: lut_data <= {-10'd04447};
        10'd 1378: lut_data <= {-10'd04378};
        10'd 1379: lut_data <= {-10'd04310};
        10'd 1380: lut_data <= {-10'd04240};
        10'd 1381: lut_data <= {-10'd04171};
        10'd 1382: lut_data <= {-10'd04102};
        10'd 1383: lut_data <= {-10'd04033};
        10'd 1384: lut_data <= {-10'd03964};
        10'd 1385: lut_data <= {-10'd03894};
        10'd 1386: lut_data <= {-10'd03825};
        10'd 1387: lut_data <= {-10'd03755};
        10'd 1388: lut_data <= {-10'd03686};
        10'd 1389: lut_data <= {-10'd03616};
        10'd 1390: lut_data <= {-10'd03546};
        10'd 1391: lut_data <= {-10'd03476};
        10'd 1392: lut_data <= {-10'd03406};
        10'd 1393: lut_data <= {-10'd03336};
        10'd 1394: lut_data <= {-10'd03266};
        10'd 1395: lut_data <= {-10'd03196};
        10'd 1396: lut_data <= {-10'd03126};
        10'd 1397: lut_data <= {-10'd03056};
        10'd 1398: lut_data <= {-10'd02986};
        10'd 1399: lut_data <= {-10'd02915};
        10'd 1400: lut_data <= {-10'd02845};
        10'd 1401: lut_data <= {-10'd02775};
        10'd 1402: lut_data <= {-10'd02704};
        10'd 1403: lut_data <= {-10'd02634};
        10'd 1404: lut_data <= {-10'd02563};
        10'd 1405: lut_data <= {-10'd02492};
        10'd 1406: lut_data <= {-10'd02422};
        10'd 1407: lut_data <= {-10'd02351};
        10'd 1408: lut_data <= {-10'd02280};
        10'd 1409: lut_data <= {-10'd02209};
        10'd 1410: lut_data <= {-10'd02139};
        10'd 1411: lut_data <= {-10'd02068};
        10'd 1412: lut_data <= {-10'd01997};
        10'd 1413: lut_data <= {-10'd01926};
        10'd 1414: lut_data <= {-10'd01855};
        10'd 1415: lut_data <= {-10'd01784};
        10'd 1416: lut_data <= {-10'd01713};
        10'd 1417: lut_data <= {-10'd01641};
        10'd 1418: lut_data <= {-10'd01570};
        10'd 1419: lut_data <= {-10'd01499};
        10'd 1420: lut_data <= {-10'd01428};
        10'd 1421: lut_data <= {-10'd01357};
        10'd 1422: lut_data <= {-10'd01285};
        10'd 1423: lut_data <= {-10'd01214};
        10'd 1424: lut_data <= {-10'd01143};
        10'd 1425: lut_data <= {-10'd01072};
        10'd 1426: lut_data <= {-10'd01000};
        10'd 1427: lut_data <= {-10'd00929};
        10'd 1428: lut_data <= {-10'd00857};
        10'd 1429: lut_data <= {-10'd00786};
        10'd 1430: lut_data <= {-10'd00715};
        10'd 1431: lut_data <= {-10'd00643};
        10'd 1432: lut_data <= {-10'd00572};
        10'd 1433: lut_data <= {-10'd00500};
        10'd 1434: lut_data <= {-10'd00429};
        10'd 1435: lut_data <= {-10'd00357};
        10'd 1436: lut_data <= {-10'd00286};
        10'd 1437: lut_data <= {-10'd00214};
        10'd 1438: lut_data <= {-10'd00143};
        10'd 1439: lut_data <= {-10'd00071};
        10'd 1440: lut_data <= {10'd00000};
        default: lut_data <= {10'd99999};
    endcase
end
endmodule
